ELF              d  4   �.      4    (                 �  �           (  (  (  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �z    ��   ��t���   ��t��1�ÐS���V  ���  ��������Q�������[Ív WVS�3  ���  �|$��   ��t9���   ��t/�Љ��gfff���������)�t������   ���   9�r�[^_Ív 1ۅ����ڍv VSQ��   ��\  ��   ��t&��j�S�Ã���t��   ���   ��C   ��Z[^�S���~     �\$��   ��t��t���   +������[Ð1���[ÐS���B   �  �\$��   ��t��t���   ���[Ív �   �  �T$��   ������Ë$Ë$Ë4$�                                                        	4D  �         �W�������� ��Bw ����timer                                 @                      ticks                               seconds                         $   sleep                           L   sw_new                          �   sw_ms                           �   sw_rst                          4  (                        �  ���o�     0     �  
   k            �     8               ���o                                                           S   4  -     b   d       #   L   e        $   %     ?   �   ;            #     /   �   D      timer_get_ticks timer_get_seconds timer_sleep timer_sw_create timer_sw_elapsed_ms timer_sw_reset cdl_main  (     `     �     �     �     �                 �  4                   2   �  ^   E   D  	S   X   r   r   r   r   r    int �  
�   �   �   r    =  �   �   �   r   r   r      �   �   �   r   r    0   X       �  #       	2    O      ,  	2     	^  �   
^     4n    	r   �   n  	2    �   ~  	2        ,  �	E  �  U   /  p  �  �  �   �    �     �  �  !�  �   "�  �  %   �  &  $H  '"  (�  (;  ,�   )�  0�   *�  48   +�  8k   .h  <�  /�  @a  0�  D�  1�  H�  2�  L�  3  Pk  46  T�   5Z  X6  8t  \�   9�  `d  :�  d   ;�  hA  <�  l�   =�  p�  >�  tQ  ?  x�   @�  |�  A-  �T  BA  �-  CV  �e  F`  �X  G`  �#  H`  �}  I  �#  J`  �    M  ��   N�  ��  O�  �k  P�  �  Q�  �3   R  �[  S8  �x  T[  �   Uo  �  V�  �2  W  �H  X  �P  [�  � P  P     E  E   i  i   �  Z  E   �  E   i   u  �  E    �  �  r   �  P   �  r   �  P  P   �  �  �  r      �  r     P  �  r    �  r   "  P  E   r    	  r   ;  P  r    '  9   h  P  r   r   G   y   �    @  �  r   r   r   r   r    m  �  r   r   P  r    �  �  r   r   P  r   r    �  �  r   r   P   �    r   r   r   r   P   �  6  r   r   r   r   r   r      U  9   U  r   �    ~  ;  t  E   r   i   _  �  E   �  i   �  y  �  �  P   �  �  �  P  i   �  r   �  P  P  i   �  �  �  P  r    �  �    P  P   �  r   -  �  P     i  A  P   2  V  r   �   F  &   [  z  z  z  z   r   e  r   �  r   r   r    �  r   �  r   �  r    �  r   �  r   �  i  r   �  r    �  r     r   �  i  r    �  r   8  r   E   i  r   E   z     r   [  r   E   i  r    =  r   o  r    `  r   �  �  �  �   t  �   ]�  $_	�  �   _   �  _'E        _3�  ,`		  �   `   +   `)r    �   `6r   $�   `R	  ( �  y   `]�  	  �  sys "	  $  (	]	  �  )&    }  *	r    5  +9	  �  y	  	2    �   Gi	  @  �  P	     �  W	  d     ��	  api W'"	  �  I   A4  -   ��	    AE   � 
sw C�	         ]	  �  7r   �   ;   �^
    7E   � 
sw 9�	        
now :&   ,   *   s  ;&   8   4    o  -E   �   D   ��
  
sw /�	  Q   M    �  L   e   ��
  ms r   � >  &   f   `   �  &   �   y   B   &   �   �      r   $   %   �  8       _  

&       #   �  I   :;9I8   !I  'I  '   :;9I  :;9  I  	! I/  
4 :!;9I�B  4 :!;9!I�B  $ >  4 :!;9I   :!;9I  .?:!;9!'@|   :!;9I  %     $ >  & I  :;9   '  &       'I  4 :;9I  .?:;9'I@z  .?:;9'I@|  .?:;9I@|  .?:;9I@z  H }   . ?:;9I@   �          ��S    ��S���    ��P    ��p s ���P     ��P��S       v{P{�Q��Q         ��s p ���S��S��r 3&p �   ��S                            �    7   �          D   L   <   <   ^        	�f J f J& 0M� X��!	f J fLK3X�.01	= �M xt .��fK%�	uf f	/w'h!f JKg1<=J  y.5#h!f JK f/,��	� g ping close strncpy cdl_symbol_t menu_def_t version send fs_exists target timer_sw_reset label win_handle_t create_window cdl_exports_t my_symbols socket memcpy strncmp lib_name symbol_count set_window_menu memmove fs_delete fs_rename free get_launch_args kernel_api_t sendto exec net_get_interface_info malloc memset mouse_cb_t fs_list process_events timer_get_ticks timer_sw_create exit timer_sleep fs_create draw_image_scaled draw_image input_cb_t draw_text_clipped my_exports sprintf strchr cdl_main fs_read print uint32_t item_count menu_cb_t mem_total itoa dns_resolve start paint_cb_t char strlen recvfrom strcpy draw_rect_rounded get_kbd_state realloc action_id timer_sw_elapsed_ms GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection exec_with_args func_ptr long unsigned int draw_rect timer_get_seconds items handle get_fs_generation stopwatch_t strcmp http_get strstr mem_used draw_text connect diff recv running ticks_to_wait fs_write bind start_tick /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/lib/timer.c usr/lib usr/lib/../../sys cdl_defs.h       ���� |�             #          $   %   A�C_A� ,       L   e   A�A�A�S
�A�A�D 0       �   D   A�A�AXB H\A�A�   (       �   ;   A�Cm
A�BEA�          4  -   A�CgA�        d                        �            �                                 ��	   $             ,        @  �                  ��#   �        9   (        B           X   �        n           �   $   %     �   �   ;     �   4  -     �       #     �   L   e     �   �   D     �   d        timer.c sys my_exports my_symbols __x86.get_pc_thunk.si _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ timer_get_seconds timer_sw_elapsed_ms timer_sw_reset timer_get_ticks timer_sleep timer_sw_create cdl_main  .symtab .strtab .shstrtab .text .gnu.hash .data .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                         �                 %         �  �  4                !   ���o   �  �  @                +                                 1                              :         $  $                    ?         (  (  �   	             H         �  �  �   	            P         0  0  k                  X              �                   d              �  �                 r              �!  �                  �              �"                     �              �"  �                 �      0       t$  �                �      0        *  i                 �              �*  4                 �   	      �  �  8                              �+                 	              �,  �                                �-  �                  