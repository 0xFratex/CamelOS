ELF              �  4   �6      4    (                 
  
           �  �  �  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      UWVS��8�  ��  �D$L�D$�L$P�T$T�T$ �t$X�t$$h�VRQ�L$8��P���  �P@����
�D$,��,   �L$<�q
��v  �� ����Ɛ�; th � �SU�t$���  �QD����-��9�uڋL$�D$���h000�j�t$(�D�P�t$,���  �P@���  �D$l�����������T$h���\$d�T$,�T$`�@D��L[^_]��UWVS���  ��  �|$0��   �D$� ����   ������,   �L$Rj-j �L$�P���  �P\�������   �\$�+��    �)��\� �D$�1�����,t�@���u��)��T� �L$�� E�D$�(��������P���  ��<$���  ����  �������T$@� ��,[^_]����,   �D$�Í�I  �|$f���Pj-j S���  �R\��-XZSW���  �Pd��9�u؋|$Qj-j �D$I  P���  �P\�D$�    ���I  ������D$�(1���    �%����WVS��t�  �é  �|$ W�t$V������P���  ���   ����u_��������P�L�����V������P�t$<V���  ���   �4$�(�����W������PV���  ���   �4$��������p[^_�f���������P���������p[^_Ív VS��   �i  ���  ��$�   ��߃�L��   ��Wti��P��   ����'���P������j@�t$V��:���P���  ���   ���xjPV��B���P�t$LV���  ���   �4$�X������Ą   [^Ã�������P�=���������$�/������Ą   [^Ív �����Ą   [^�f�����L���P�������Ą   [^ÐWVS�   ��  �D$���  ��,   ��v  �f����  Qj-j S�P\��-��9�u����_���P������XZj ������������h�   h@  ��t���P���  �P<�� �����1�[^_Ë$Ë4$Ë<$�  Keys: [L] List [P] Ping [W] Wifi [NetTools]  
 eth0 1. eth0 (RTL8139) - UP    IP: %s    MAC: %s No active interfaces found. [WIFI] Scanning... No wireless extensions. Pinging 8.8.8.8... 8.8.8.8 Reply: %s Request Timed Out. NetTools v1.2 Ready. Network Tools                                                           a0!         ���0��a����	�|��8�.m�G      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �  ���o�     �	     D	  
   E            
                    ���o                                                           &   `  �     <   �  �     
   @  v    3     �            �                   �   o     on_paint log_buffer net_log log_head cmd_list_dev on_input cdl_main              �       y             �      �  1   �  P   C     	P   U   o   o   o   o   o    int �  
�   �   �   o    -  �   �   �   o   o   o    �  �   �   �   o   o    0�   J   �    o  #   	    1        	  #  1     	R  �   
R   �  4b  �  	o   � 	  b  1    	�   r  1        #  �	  �       -  g  F  �   V  Z  \     p  �  !�  �   "�  �  %�   6  &�  $8  '�  (_  (�  ,�   )p  0�   *�  48   +p  8]   .%  <�  /I  @  0h  D�  1�  H{  2�  Li  3�  P1  4�  T�   5  X&  81  \�   9Q  `*  :f  d   ;�  h�  <�  l�   =�  p�  >�  t  ?�  x�   @Q  |�  A�  �  B�  ��  C  ��  F  �  G  ��  H  �Y  I<  ��  J  �    M�  �y   NZ  �?  Ox  �   Px  ��   Q�  �3   R�  �!  S�  �(  T  �   U,  �  VJ  ��  W�  ��  X�  �@  [\  �          C   &  &   �    C   F  C   &   2  V  C    K  [  o   p     a  o   �       u  �  �  o      �  o   �    �  o    �  o   �    C   o    �  o   �    o    �  8   %    o   o   E   v   �    �  I  o   o   o   o   o    *  h  o   o     o    N  �  o   o     o   o    m  �  o   o      �  �  o   o   o   o      �  �  o   o   o   o   o   o    �    8     o   �    r  �  1  C   o   &     K  C   K  &   P  6  f  �     V  �  �    &   k  o   �      &   �  �  �    o    �  �  �       �  o   �  �     �  &  �     �    o   �     &     7  7  7  7   o   "  o   Z  o   o   o    A  o   x  o   K  o    _  o   �  o   K  &  o   K  o    }  o   �  o   K  &  o    �  o   �  o   C   &  o   C   7   �  o     o   C   &  o    �  o   ,  o      o   J  �  �  �   1  �   ]}  $_	{  �   _   �  _'C        _3Z  ,`	�  �   `   +   `)o    �   `6o   $  `R�  ( {  k   `]�  �  O  sys �  �  	   	  1   1   , O  �  @  P  	o      �  H�  �  �   ��	  api H'�  � 
win LC     )   u	  i Jo          N  �
  �  [
    �   7�	  !key 7o   
buf ?�	  
res Ao   
msg C�	     	  �	  1   ? -  +    �   �[
  x +o         y +o   #   !   w +!o   -   +   h +(o   7   5   "B   -	o   E   ?   #   i .o   b   `     $C  `  �   ��
  ip  
�   ��mac  �
  ���  S   �
  buf #�	  ���  �
  �  �
  �  �
     �
   	  �
  1    �  �   o  �,  msg   m   i   i 	o   �   ~   %�  (   
i o     &�	    �   �'�	  � (�	  D      7�  )�	  �   �   *�	     �	  ��~+�	  �   �   ,�	  v  "   �  �	  ���  �
   S  �
  �  �
    �  �
  �  �
  �  [
     I   :!;9I8   !I  'I  '  H }   :!;9I  ! I/  	I  
4 :!;9I   :!;9I�B  :!;9  4 :!;9I  $ >  4 :!;9I�B  4 :!;9I?      .?:!;9!'@  4 1  %     $ >  & I  :;9   '  &       'I  .?:;9'I@|   :;9I   .?:;9'   ! :;9I  "4 :;9I�B  #U  $.?:;9@|  %  &.1@|  ' 1  (1R�BUXYW  ) 1�B  *1U  +4 1�B  ,1   �          ��0�    ��     ��    ��    ��      F\�\#
�\kVk��\#
�  Fk0�     ��� ���       ��0���P��0�    ��� ���     ��P��P                  �          &         FUl� ���� ���� �    7   �         L   U   	   	   h   +     *.u	 	�t�Y  d �Jt�f��t�=sW.Y��Xf�.�	� Y	Y!	=
<NKu   1 �4 1 f �/1 s .rt#.�& � 	xJun	a
�	 �	u�- �	�/ t�	�"�//]y�	�	�g@ ��	t���	
<# r�Y���,�!	g	 ' �$ f  � �*� ping close strncpy cdl_symbol_t menu_def_t version send fs_exists start_y label win_handle_t create_window cdl_exports_t socket memcpy strncmp lib_name symbol_count set_window_menu on_input memmove fs_delete fs_rename free get_launch_args kernel_api_t sendto exec net_get_interface_info malloc memset mouse_cb_t fs_list process_events log_buffer exit fs_create draw_image_scaled draw_image input_cb_t draw_text_clipped sprintf strchr cdl_main fs_read print uint32_t item_count menu_cb_t mem_total itoa dns_resolve paint_cb_t char symbols strlen recvfrom strcpy draw_rect_rounded cmd_list_dev log_head get_kbd_state realloc action_id GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection exec_with_args func_ptr long unsigned int draw_rect get_ticks items get_fs_generation strcmp net_log http_get strstr mem_used draw_text connect recv on_paint fs_write bind usr/apps/nettools_cdl.c /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/apps usr/apps/../../sys cdl_defs.h      ���� |�  l           �   A�A�A�A�CLlPATAXA\G`h@QDAHALDPL@XLEPBTDXE\D`vA�A�A�A�   �       �   o  A�A�A�A�C0y4B8B<G@N0Z<G@hA�A�A�A�B0����[4B8B<A@M<A8A<A@L0I4B8B<J@V0   �       `  �   A�A�A�C�P�E�G�O�G�G�H�A�G�E�W�A�G�A�W�C
A�A�A�CC�G�H�CA�A�A��         �   A�A�F�o�G�H�B�E�G�N�E�A�G�E�W�F
A�A�AC�G�V�F
A�A�DK
A�A�CC�G�H�FA�A� X       �  �   A�A�A�lBBA IGG HABF F$E(E,G0LH�A�A�        �            �            �                                 ��   �                    ��   �        *   �        @   �        I   �        _           u   `  �     �           �     �     �       �     �   �  �     �   �   o    �   @  v     nettools_cdl.c sys __x86.get_pc_thunk.si __x86.get_pc_thunk.di _DYNAMIC __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ cmd_list_dev log_head on_input on_paint cdl_main net_log log_buffer  .symtab .strtab .shstrtab .text .rodata .gnu.hash .got .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_rnglists .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                           �                 !      2   �  �                  -         �  �  4   	             )   ���o   �  �  @   	             3                              8                              A               �                  F         �  �  �   
             O         D	  D  �   
            W         �	  �  E                  _                �                 k              �%  R                 y              G(  �                  �              )                     �              +)  *                  �              U)  �                 �      0       �+  D                �      0       1  s                 �              �1  �                 �   	      
       	                           T4        	         	              T5  �                                6  �                  