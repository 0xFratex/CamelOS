ELF              Lz  4   �9     4    (                 �� ��          �� �� �� �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      WVS��� ��u/�Nf��p����w�� �q����w�� 8�uG�J���t���
��u�)�[^_�����)�[^_��J1����
1��ߐUWVS��<�3�  ��(�  �ŉЅ�t
��|  ��t,�������0   ���   �   ��6�J  ��(����㐍������0   ����܍v �D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   ��   �D$    �D$    �D$    �$�  �   ������   ��} �u�]�<$�}�|$�}�\$�]�t$�u�U�M �T$�U$�|$�}(�\$�]0�T$�U4�t$ �u8�|$$�}<�L$(�M@�\$,�]D�T$0���   ���   ���   �D$4���   �D$8���   ���<[^_]Ív �L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �������L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �   �}����L$�D$8   �D$4    �   �D$0�����D$,    �D$(   �D$$   �D$    �D$   �D$   �D$    1������D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$   �D$    �D$   �D$   �D$    �D$    1������v �L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    1��D$    �D$    �D$   �$�  �   ������   ��\�����D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$    �D$    �D$    �D$    �D$   �   ������L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    1��D$    �D$    �D$    �$�  �   ������   ��l�����D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   �   �D$    �D$    �D$    �$�  �   ������   ��������L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$   �D$    �D$   �D$   �D$    1��D$    �D$    �D$    �$�  �   ������   ��H�����D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$
   �   �   �D$    �D$    �D$    �$�  �   ������   �������L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$   �D$    �D$   �D$   �D$    1��$����v �L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �������D$8   �D$4    �   �D$0�����D$,    �D$(   �D$$    �D$     ����f��D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$   �D$   �O�����L$�D$8   �D$4    1��D$0   ��D$,    �D$(   �D$$   �D$    �D$   �D$   �D$    1��D$    �D$    �D$    �$�  �   ��f �������������D$8   �D$4    1��D$0   ��D$,    �D$(   �D$$   �D$    �D$   �D$   �D$    �D$   �   �   �D$    �D$    �D$    �$�  �   ������   ��<�����L$�D$8   �D$4    1��D$0   ��D$,    �D$(   �D$$   �D$    �D$   �D$   �D$    1��o����v �L$�D$8   �D$4    1��D$0   ��D$,   �D$(    �D$$    �D$     �D$    �D$    �D$    1��D$    �D$   �D$    �$�  �   �������f ��P�����D$8   �D$4   1��D$0�����D$,    �D$(   �D$$    �D$    �D$   �D$   �D$   �D$   �   �   �D$    �D$    �D$    �$�  �   ������UUU�������D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$   �D$    �D$    �W�����D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$   �D$    �D$    �D$   1�������v �L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    1��D$    �D$   �h����v �D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   ������L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    1������v �D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   �(����D$8"   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   �   �D$    �D$    �D$    �$�  �   ������   ��������D$8   �D$4    �   �D$0�����D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   �)�����D$8   �D$4    1��D$0   ��D$,    �D$(    �f�����D$8   ��f��D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$   �D$    �D$    �D$    �D$    �D$   �   �   �D$    �D$    �D$    �$�  �   ������   �������L$�D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �   �D$   �D$    �D$    �$�  �   ������fff������f��D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$   �D$   �D$    �D$   �   �`����D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   �   �����v �D$8   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   �   �D$    �D$    �D$    �$�  �   ������   �������D$8(   �D$4    1��D$0   ��D$,    �D$(    �D$$    �D$     �D$    �D$    �D$    �D$   �   �   �D$    �D$    �D$    �$�  �    ������   �������UWVS���7�  ��(�  �Ë��\ =�   ��   ��  ��   �< �<$Ǎ,�����.�\ ���\ �T$�O�L$$�O�L$(�O��d  �O���  �o���  �l$�o���  �l$�o���  �o ��  �o,�_0�����   ��1ҁ�   ��<$������|$�T$�L$��~}1ɋl$�����<$Ǎ<��<��l$�L=(���  ��~)�$����\$�D(   @���\ ��[^_]Ív ���  ��͋��  ��Ë��  ���	�ũ�[^_]�f�1��1��\����UWVS�����  ����  �Ê < u	f�C�< t�<#��  ��d����������ƅ���   �S�C��u�  �v B���t<(u�B�
�A�<	�{  1����� B�A���؊
�YЀ�	v������B�
���5  ��0��	w��HЀ�	�    ��  f����	B�H���ي�XЀ�	v����  �v ��h������S�������  ��n������>������+  ��t������)������  ���������������  �����������������  ��%��������������  ��x��������������  ��}��������������  ��������������\  ��������������G  ����������������  ���������l�������  ���������W�������  ���������B������W  ���������-�������  ���������������K  ���������������J  �����������������  ����������������*  ����������������  ���������������  ���������������4  ����������������  ���������p�������  ���������[�������  ���������F�������  ���������1�������  ����������������  ���������������v  ����������������  ����������������  ���������������}  �� ������������^  ��,������������?  ��3������������   ��;������t������Q  ��B������_������2  ��I������J�������   ��[^_]�f��s����E V���   �ǃ�����   ��s	��D$1����0	�9L$t)A9�t$����ZЀ�	v�j����w ��W	�9L$uؐ���   ���[^_]�f��j����w���7	�묍v B���t.��0<	w��{Љ�<	w�v �4��B��0��ފ�C�<	v�	�	��   ��1���   ������**������1�����1�1��и������������ �������� ������������������  �������� � �����������������  ������ ����������������� � ������  ������� ���������� ��y����P���o�����  ��e����� ���[���� ����Q���������G�����ح��=����<���3����� K��)���� ���������·������r�������������������������������������������������������Gc��������S����B�<	�    w�v �����0���A��ZЀ�	v��et��pu�ytt[�f��ymu�� ����[Ð� ����9��8�������)�[Å�t�8 t념1�ÐVS�0�  ��!�  �Í�U����v�����u[^Ív ��Z������_�������   ��`������J�����tz��g������9�����tu��n������(�����t|��u�����������t_��|�����������tf���������������t_����������������������b����   [^ø   �P���f��   �D���f��   �8���f��   �,���f��   � ����   ����VS�(�  ���  �Í������n�����u
�   [^�f����������S������  ���������>������r  ���������)������I  ���������������\  ����������������S  ����������������&  ����������������5  ����������������*  ���������������  ���������������  ���������������	  ���������l�������  ���������W�������  ���������B�������  ���������-�������  ����������������  ����������������  �����������������  �����������������  �����������������  ����������������  ����������������  ����������������  ���������p������t  ���������[������U  ���������F������6  ���������1������  ����������������  ����������������  �����������������  �����������������  ��0��������������  ���������������q  ��!������������R  ��������������3  ��������t������  ��������_�������  ��������J�������  ���������5�������  �������� �������  ��"������������y  ��'�������������Z  ��.�������������;  ��5�������������  ��9�������������  ��>�������������  ��F�������������  ��N������x�������  ��T������c�������  ��[������N������b  ��f������9������C  ��n������$������$  ��v������������  ��|��������������   ������������������!�s����   �i���f��   [^ø   [^ø   �M���f��   �A���f��   �5���f��   �)����	   �����
   �����   �����   �����   ������   ������   ������   ������   ������   ������   �����   �����   �����    �����   �����8   �����7   �����6   �u����5   �k����4   �a����3   �W����2   �M����1   �C����0   �9����/   �/����.   �%����-   �����,   �����+   �����*   ������)   ������(   ������'   ������&   ������%   ������#   ������   �����   �����   �����   �����   �����   �����   �{����   �q����   �g���U��WVS��\  �b�  ��S�  ��E ���  ��j��u�u�u�u�P@��h����j�u�u�u��E �P@�E��
�������� ����������
  �E����������H0 �]1��������������������������������9�(/ ��  �������Pjjv������S��E �P@����������E ���   ����~�   ������PR��������������������E �Qh������Ƅ���� ����������~	fǅ����..h   ��������������CP��E �PD���������  hfff��������������ChP��E �PD��xG�������  ��;���������f�hfff���N���R�������CP��E �PD�$����j$�u�E��P�u��E �P@��h����j�u�E��@P�u��E �P@�E�x"�E��
��������jj�jjWP��E �PT�E�X*�� h   �������PS�E��P��E �PDXZjj�jjW�E��(P��E �PT�� h   ���^���PS�E��.P��E �PDYXjj�jjW�E��FP��E �PT�� h   �������P������S�E��LP��E �PD�E��V����E�XdXYjj�jR������WS��E �PT��h����j������RWS��E �P@�E�Hi����  �� �8 �  h   �P������Q��������E �PD����  @�   �������  ����/��h   �jj�E��&P����  ��������P��E �P@�� �E�M���������jj�jjW�D�P��E �PT�� h   �������P�������C�P��E �PD��H   ���8 t#h����P�E�}�D8�P��������E �PD���E�xD�������E)�+E���������M�Y쉝������j�PQW�u��E �P@��h����j�uW�u��E �P@��(   ������� ���������������� ���\ ����  ���\ ǅ����    ������������ȉ��������f���������������49��\ ��  �{ϋ�����)ǋ�C�������9ȉ�����|�9�����|�������������S$��t_�C ��E �R@�������S�������S����������  ��������������������������W�������������Ѓ� �������C(���:����C�������C�S�������S�{ ������������������������������PR������W��������E �P@��������������Q������R�������:)�P��������E �P@�������	������)�σ�������������RQW��������E �P@��������������������QW�������������)�P��E �P@�� �������>���f���x����������#���f�����������������   ���Ѝ�ЍG1���  9�}�Ё��  9�uꉝ�����H������9�}]����E h�����������}�   Pj��������������ȅ��  �����Й���������V��������
P�S@�� �e�[^_]�f�h����������P������Q��E �PD���%������������ ��~E��4��������� ������������É������]�K	������������1��������������5  �)ЋM�D
��  �����������  =�  �  ��y������������W��E ���   ��������9��^  PQW������������P��E �Ph������Ƅ���� ��������������S��������E �PD�����  ��t8����������E ���   Z������j��P�CP��������E �P@�� ��  �  u#������������S������@P��E �PD��f���������������� ���  9�������������  ������)Ë�   ������9�|�9�����|�������)���~���(  ��tt����  ������ȉ�����������������9������Y����������������Q�����W������������P��E �Pd������f�ǅ����    �N����������+�  �������E������냉�������� ���������������������Ћ�����)�PW�������������Q�������Ѓ�������������������)�P�������������9R��������E �R@��������������QQW��������E �R@�����������������)ʃ�������QQW������R��E �R@������������)ȃ�������QQ������P��������E �P@��������������QQ��������������E �P@�� �������s���ǅ�����   ������������E+�  ���������&����v ��������]�`���UWVS����  ���  �$�Ջ���  ���k  ����  ���U  ���M  �$�ȍ��v @9��7  �8 ~�I ��  �   �G��I ��    �D$����������(I ��T$QhD  j �D$P��E �P\�D$�    �E�$��E �P�T$��(I �B(�T$����t!RU�t$P��E �P`�T$�B(�( �j,������  ��t�D$����������`  ��`  �0   󥉐   ��$  ����   ��(  �t$��,  �D$��(  �zu'��~�   P��E U�t$���   S�Ph�+ ����[^_]Ë���  ����  �WU�t$����  P��E �P`���  ����[^_]ËD$��$  �y���UWVS��  �D�  ��5�  �ÉT$� �l$?����   �v < ��   �P�����   ����   1����?��   CB�D �����   <:u��D@ C��< t<	uC��v 1ҍL$��u�   ���twCB����tl<;u�Ƅ�    C�|$@���������������uV��$�    �X  ��$�   �����|$�����@�����  [^_]ÐC��,����D@ �f���f�Ƅ�    �f���������������uY��$�    �2  ��$�   �-����|$�G�Ƅ$�    �|$@���������G�������   ���������2�������   ��������������t���������������uG��$�    t-��$�   ������|$�G��~��H�����GH   �����D$�@   �������������������u6��$�   ����������������   �D$�@�  �����   ��������������m�����u0��$�   �������W����������|$�G�y����   ���������������,�����uW�������P��$�   P��E �Px���������|$�G�,�������������������M����D$�@�  ������������������u(��$�   ��U�����������uQ�D$�@   �������,������������D$ul��$�   ��7������o������L$u1�D$�@ ����������&������J�����up�D$�@   �l�����$�    t	���������D$�H �M�����<������
������D$ul��$�   ��7�������������L$u1�D$�@$����������������������up�D$�@   �������$�    t	���������D$�H$�������J������������D$ul��$�   ��7������m������L$u1�D$�@(����������������H���������|$�G�j�����$�    t	���������D$�H(�K�����V������������D$u0��$�   ��7�������������L$�q  �D$�@,����������c�����������D$����  ��j�����������u"��$�    t��$�   �����|$�G0������v������w�����u"��$�    t��$�   �M����|$�G4�������������D�����u"��$�    t��$�   �����|$�G8�T�����������������u"��$�    t��$�   ������|$�G<�!��������������������   ���������������u"��$�    t��$�   �����|$�G@�������������������u=��$�    t��$�   �j����|$���   ���   ���   ���   ���   �������������F�����ul��$�   �����|$���   �]����|$0�|$�   󫍼$�   �? ��  ��u��   G�? t�B�T$���L����L$�T$�D���G��u��ō��������������u,��$�    t��$�   �s����|$���   ������   ��ꍖ��������������  ���������w������N  ��$�    �	  ��$�   �E����|$���   ���y���Ǉ�      �j������a����D$0�|$�G0�D$4�G<�D$8�G4�D$<�G8�<����|$ �|$�   �|$0�|$�   󫍼$�   ��7����D$�����   �|$��   < uG�? t��T$����������   �L$�T$��   �T$�L$��A�L$���u�f�G���t�< u�똀�$�    t	���N������D$�H,�����|$��   �|$�p�������|$0 u�D$ �|$�G ����|$4 u�D$$�|$�G,����|$8 u�D$(�|$�G$����|$< u�D$,�|$�G(�����|$u�����|$0 u�D$ �|$�G,�G(�G$�G �������������������|$0 u�D$ �|$�G$�G ����|$4 u�D$$�|$�G,�G(������u*�D$0�|$�G<�G8�G4�G0�����D$1ɉ��   �}������
����D$0�|$�G4�G0�D$4�G<�G8�W�����������������u~��$�    tc��$�   ������|$���   �������������$�   �? uG�����-����L$���   ���   ���   ���   ���   ��tRG���D$1҉��   �������������������uF��$�    t+��$�   �[����|$���   �����������? uRG���D$1����   �q�����
������.�����uW��$�    t<��$�   �����|$���   ��������3������f����L$���   ��tbG���D$1ɉ��   �	�����������������uY��$�    t<��$�   �����|$���   ��~!��0�����Ǉ�   0   �����< uOG���D$ǀ�      ������"������\�����ua��$�   ��-������D�����u$�D$�@   �f������^�����������m�������������������   �D$�@   �-�����<�����������D$��uz��$�   ��E������������t;��M�����������tG��T�����������t,��7�����������u�D$   �D$�|$���   �����D$   ���D$   �ٍ�[������[�����up��$�   ��M������C�����u4�D$ǀ�      �b�����4���������������|$�G�A�����f����������������|$���   ������o��������������   ��$�   ��x�����������tZ������������¸   ��tB���������������S  ���������������4  ���������k������������|$���   �������������D�����u%��$�    t��$�   �����|$���   �Q����������������D$��uk��$�   ��o������������tC�����������������  ����������������f  ��������������u�D$   �D$�|$�xL������������������D$����   ��$�   ���������n�����tm���������]�������  ��-������H�������  ���������3������  ��	�������������  ��������	�����u�D$   �D$�|$�xP�#�����#��������������   ��$�   ��/����������������   �������������   ��to�L$���������������L$tV���������~������P  ���������i������;  ��-������T������  ��7������?���1Ʌ������D$�HT�_�����@����������D$����   ��$�   ��7��������������   ����������������  �����������������  ����������������  ����������������  ��-�������������  ��/������~�������  ��7������i�����u�D$   �D$�|$�xX������K������@�����uS��$�   ��U������(�����t/��P����������¸   ��t��\������������������|$�G\������i������������u"��$�    t��$�   �����|$�G`�������s�����������u"��$�    t��$�   �����|$�Gd������������v������D$uK��$�   ��7������Z������L$t��$�    t	���1������D$�Hh�i����D$�@h�����Y������������������   ��$�   ��U������������uL�D$1҉P`�Pd�@h���������D$   �t����D$   �g����D$   �Z����D$   �M�����7����D$��藿�����A  �D$�@`   �@d   �@h�����������������d�����u"��$�    t��$�   �:����|$�Gl�t������������1�����u"��$�    t��$�   �����|$�Gp�A�����������������u"��$�    t��$�   ������|$�Gt�������������˾����u"��$�    t��$�   �����|$�Gx�������������蘾����u"��$�    t��$�   �n����|$�G|�������������e������������$�   �? uG���? uG���������L$���   ��t"G���������L$�A`����K���< tG��? u#G��G���^����L$�Ad����#���< tG����?����L$���   ��t*G��G�T$���������������������|$�Gh������? uG���D$   �����D$   ������������L$���   ��t_G���D$   �a����D$   �����D$   �����   ������   ������   ������   ������D$   �����< uG�����4����������|$���   ����UWVS��   �$ ��<  �n�  g�  �D$����   �  �D$����  ���������WR�D$��E �Px������  �P�< ��  �H�����  <(u�f�B�< t��H���v�<"t<'u��r�t$ �R1ɍ�$/  ��tM�ŋ\$ �f�C����t5��8�t/���  t'A��\u�C��t�<n��  ��  ������uˉ\$ Ƅ0   ��$0   �L  ����$<  U�\$��E ���   �Ɖڍ�  ������~�  �  ��U�����P��E �Pd3��$@  ������  ��$/  �t$L�l$�|$8��t$�FF�t$����  <<��  < ~��D$� ����  �\$��C���t<<u��ދD$)ƅ���  �D$�
�v N�  �|0� ~�D$��I ��  �b  �B�L$��I ��    �D$Ѝ���ЉT$$�<�    ��(I �D$�,PhD  j U�L$��E �P\�E    �F�$�L$��E �P�L$��9(I �|$(�G(�����T$$��   �T$$WV�t$P�|$��E �P`�L$(�A(�0 �q,��`  ���������0   ��󥋂��  �����T$$��   ���  ��t�t$ǆ�     ǅ`  �  ��L$э���ыt$���   ��$  ����  ��(  ��,  ��(  ��\$�L����B������<  [^_]Ë|$8�T$ �������\$�"���<r�:  <t�j����	�c����D$�@</�U  �D$�T$1���B�< t�<	t��T$1ҍ�$  ����   �\$�CB������   <>t< t	<	t��u��\$�Ƅ   ����  1ۋL$�|$L����  tAC����t<>u�Ƅ0   A�L$��L$Ƅ0   �D$��E ��u'����   �D$� �4���Ƅ$   Ƅ$0   ��t�D$����  ��tӋ�   ��tɍ�$  ���������  �D$����  먰
�8�����1����\$Ƅ   Ƅ$0   �D$��E ��u�1ۍ�$  ���x������@ԃ��Z����L$0��*�M����l$��I �L$(��  �3����A��I ��    �D$H����D$D��������(I �T$�D$�RhD  j �D$0P�W\�T$4�   �=(I �|$D�D$,�|$@��,I ��jV�t$ �D0P��E �Ph�t$`����  ����蘷���T$4��`  �0   󥊄$@  ������  ��$0  ��0  �t$@9��p  �t$�\$�t0�t$<�Ή�< ��  �P�����  ���@  ��<=��  <>t< tF���u��)؉D$�  ��$0  �@   1����D$���������}�����u�|$�  �D$���������]������M  �|$�o  �D$���������9����D$��]������(�����u�|$�Z  �D$��������������u�|$�9  �D$��������������u�|$�1  �D$���������ȵ����u�|$�h  �D$��������訵����u�|$��  ���t�\$@9�������D$����  ��tA�T$H�t$(�����t$���   ��$  ����  ��(  �t$$��,  ��(  �t$0��w� ����������D$�t$$����  �s����v C������t$�F����   ������$  ��(  ��\$�z�����)؉D$�>�����$0  �@   1����F<"��  <'�x  F����u����<>tG���t< u��)��P����   wRPVU�D$��E �Ph���������Ph�   U�t$H�\$��E �Ph�D$T�|$8��������\$DǄ�     �\$$Ǆ`  �  ����o����|$���������������������|$�����PjU�D$(�\$ ��0  P��E �Ph���&���Pj?U�D$(�\$ ���  P�D$��E �Ph��������t$$��$  ��(  �I���1���Ӄ~t9��   �މ\$,���u�D$����  �D$����  ��   �������������tߋD$�t$,����  �ύN�V�΄�u�0f�F���t8�u���)ȍP����   wWPQU�D$��E �Ph���> �S���F�M���Ph�   U�D$(�\$ ��0  ����Pj?U�D$(�\$ ���  �����WjU�D$(�\$ ��0  P�\$��E �Ph���������z������������iD$(D  ؋\$4Ǆ�     ����Sh�   U�\$(�|$ ��;@  P�D$��E �Ph����$0   �������;`  ���b����p���QjU�D$(�\$ ��@  �E���Ƅ$0   1��4���f�WVS胉  ��p�  ���C�����*tN����  ��0����  ��u��C��覱����tB��   ��t�;t�[^_Ív ��+u�Ǉ��      [^_Ð����  ��u����  ��~�[^_Ë�   ����  [^_�Ǉ��      ����  Ƅ��   �K���Ǉ��      딍v UWVS��  ���  �ǭ�  �|$�ÉՉL$�v�����*��  ��+�G  �@ԉT$����  �t$��I �|$4��  ��  �G��I ��    �L$8�9������<�    �|$ ��(I �D$�RhD  j �D$(P��E �P\�D$,�    �(I �T$L�T$��>,I ��jS�L$$�D9P��E �Ph����  �t$P�ًT$�T$ ��膰���D$,��`  �0   �D$�D$��9ŋT$��  �D$�L$ ��0  �t$,��0  �t$(�D0�D$$�D$�������L$�������D$�T$0f���f��< ��  �P�����  ���/  ��<=��  <>t< tE�E ��u��)؉D$�  ��$   �@   1����T$���M�����u�|$�*  �T$���3�������  �|$�8  �D$�������������D$��]������������u�|$��  �D$���������ޮ����u�|$��  �D$��������辮����u�|$�%  �D$��������螮����u�|$�g  �D$���������~�����u�|$��  �D$9�������T$0�D$����  ��tA�D$8�L$4ȍ���ȋL$���   ��$  ���n  ��(  �L$��,  ��(  ���  � �����  ��  [^_]Ív C�2���f���)؉D$�o�����$   �@   1����E<"��   <'��   �U�Մ�u�G����v <>tE�E ��t< u���)ЍH����   �!���QPRV�D$��E �Ph�������|$���������O������8����|$�-���PjV�t$8��E �Ph���D$9��h��������v Ph�   V�t$0�D$��E �Ph���D$9��9�������Ph�   V�t$4�D$��E �Ph���D$9������Y����M�U�̈́�u�S����v E�U ��t8�u��)ȍP����   ��   WPQV�D$��E �Ph�E ��<�������Pj?V�D$$�L$,���  P�D$��E �Ph���D$9������������v �D$ǀ��     ǀ��      ƀ��   ��  [^_]�Wj?V�D$$�L$,���  뜊E �w����D$�t$����  ��  [^_]�RjV�D$$�L$,��@  �c����D$��$  ��(  �����D$ǀ��     ��  [^_]�SjV�D$$�L$,��0  P�|$��E �Ph���������\�������������D$8�t$4���������t$<Ǆ�     ����Qh�   V�|$$�\$,��@  P�D$��E �Ph����$    �������`  ���9����q���UWVS��   �$ ��\  �j�  ��_�  ǃ��      ��I ����  ǃ��      ��(  ���tg1�1�1�1�L$���w+����������~��$P  �������1�ǃ��     f��FF��t����  ���V<>�9  ��F��u���V  ��\  [^_]Ív <>��  �V��>ӈD<��G벍v < �  �P����   <>��  �V</ù�>uǍF�D$�D< �O  �v �V<-u���-�{����~>��  F�X����V<!��   </��   ����߃�A����   ǃ��     �D$���D$    �   ����f�<<������V���  ������,P  ��E�����f�<>��   �V</��   �L$���  ������DP��A�L$�����ǃ��      �������v �D< ǃ��     �F�������$P  ���F�����\  [^_]Ív ǃ��     ��1��T������-��   ǃ��     ���9���f���>�^����F�D$�T$P�D$�L$�D$�C����D$�~���ǃ��      �F�t$������D< �T$P�D$�L$����ǃ��      �F������D< �D$�2���ǃ��      �F�����~-t'ǃ��     F�-����ǃ��      �F���~���ǃ��     �F���i���f�UWVS��l  �\  ��E�  ��E ����  ����$�  ����  V�Pd�4$��E ���   ����  ���8 �D$L�Ǎ�`  ����E ����  ��t����$�  W�Pl������  ��E �ǌ  9�u͉D$�������P��H   �D$\P�D$�Pd��h��  j ��(  S��E �P\��  �D$X�     ���   �D$<�  ǅI    ��hD  j ��(I V��E �P\ǅ(I     ��I ǅ�     ǅ�\     ǅ(�      ��(   �     ��h�  S��$�  ��E ���   �����
  �L$H��D$,�  �S���ǅ�     ǅ�\     ǅ(�      ��I ��$  ����  �D$   �D$T    �D$X    �D$D    �D$4    �D$8    �D$    �D$    �D$    ��E �D$��� �D$�$�v H��  ��$  ���   �Ë�E �D$���u؋C(�$����  ���t$�D$���   �D$���  �L$��h  �F��9��F�D$���t$��E ���   ����������|$���=�  ~�D$9���  �L$���O���1�1�1ҍ� �D$$�\$���9T$�v  G9\$�  �$���C< ޅ���  ��� ���  ��  ��E �B��� �|$(���   ~�D$(�   ��    �D$ Ѝ�ЉT$0��D$LR�t$,�T$�V�T$(�ƍP�Qh�D$8��T$,� �D$ ��h  ����������ǉ��D$P�.�t$4��  �|$�9��=�  �T$0~�D$9��e  �D$ Ѝ������D$�L$(�<�|$0�D$�t$��t$��  �L$8ȉ�   �D$(�L$$��L$(�D$4�L$���  �L$(��  ��  ��`  �0   ���L$(�D$��  ���  �t$��x  u�  �L$@)ȉ�������t$0��   �D$��   ��E ��t
���  �D$ Ѝ�ЋL$ǄA�      �D$ Ѝ�ЍDE �|$$��  �t$�D�D$�$�D�<
��   ��1�9\$������\$��$  ��� �����,  ����������,  ���������   ���0  �;uߋ�|  ���J�e  ���  T$�C����w��D$T    �f��L$L$�ދD$�D$1��J����v ���  ��~D$���  �L$��h  �P9����D$��|  ���H�x  �C����  ���  ���2
  ���8  ��� ���  �  �A��� �� �D$�<(�4�    �����ȉL$$�G[��0  ��R�T$0�D$���   �D$�����T$ �L$$~�$   ΍��ȍ4 �7�D$P�t$R�D7P��E �PhXZ������P�|$�D$�DP��E �Pd�L$(�T$���   �L$ �ʋt$$��  �|$��  ��`  �0   ���ǂ  �����|$Ǉ�      �D$��   ��  �D$���  �C�D$d������  �L$L$�D$�D$�����v ���������� ���  ������������E �D$�D$,�8 �x  �D$H�8��,: ����������1Ґ�H���e  �9�s�Ή�B�  ��u�����  �É����������$�  �D$H�4V�T$�RdXZ�t$4�D$H��   P��E �Pd���  ��E ���   ���8 ���  ǀ�     ���8 ����@���8 ����  ��@����  ������@%  ���  ����������$�  ��������  ��P��E �PdY^�|$4W�������������   P��E �Pd��������E ���   �������(�  XZ��$�  ��(/ �Љ���Ѝ�H/ ��P��E �PdY^��E W��(/ �	ȉ���ȍ��   P�Rd���D$P�  1���l  [^_]ËD$�T$9�}�L$L$�D$���  ���  ����  ���  �|$ǉ��D$8    �t$D���T$�T�`����   F�t$D���  �D$���  �D$4D$�C�������D$T   �D$X    �$������,  ���/����D$,�8 �������������P�t$8�D$�Pd����E �D$�a���f��L$L$�D$�����v �T$T$�D$�_����v H���@����f�1��e�����D$T   �D$X    �����v ���  �����  ����  ����  �=�  ��  ��  )�)ȉD$8���������  �t$΋|$D���L  ��   ��t	�:��  �D$4    �D$    ��  ��t$H�W����D$�T$9��G����t$�L$�D$�4����v �0 �f����t$ ��ʍ�щT$0�4	�T$�2�L$@ǁ�     ���  �T$$։��  �O0���L$0Q�T$(�L$X��
�  Q�Pd��(�  ����_�T$0�����T$\�H��(�  �H�  �T$0�L �ʍ���������T$L��ȉD$@��   �T$@��)�H�  Ћ�  �P��  �p�t$�p���  �T$@��  ���t$0�D$X�DP��E �Pd���T$\�q�������   W���   S��E �Pd��  �     ��(  �  ǅ�     ǅ�\     ǅ(�      XZ��$�  V��E �PdY^��$�  ��(/ �Љ���Ѝ�H/ ��P��E �Pd_XS��(/ �Љ���Ѝ��   P��E �Pd����H   �D$P�"�����	��   �L$�t$�$��� =�  ��   �P��� ��������R���Ѝ�Ѝ4 ��5� ��P��E �Pd���L$(��   ���t$��  �|$  ��`  �0   ���ǂ�      ǂ  @  �|$���  �C���t$�T$$���L$�L$���k  ��� =�  ��   �D$Z�����v ����D$�D$�D$������v �D$d�����f���H�D$D�|�`����   ����)��Ph�  ����躪����|  ���|����B�=�  w.��  )����D$8�������  �L$���  �T$4�j����v �D$8    1��������P��� ��������R���Ѝ�Ѝ4 ��5� W��E �Pd�L$(�D$ȉ�   ���t$$��  �|$��  �ύ�`  �0   �ǂ�      ǂ  P   �|$���  �t$$�N��P�X^�GPjT���Ʃ���C�D$Z������������ =�  ��   �P��� ��������R���Ѝ�Ѝ4 ��5� W��E �Pd�D$(�T$Љ�   ���L$$��  �|$��  ����`  �0   �ǂ�      ǂ  F   �t$���  �L$$���P�_X�FPjN���������D$P�����f��Ӆ�������=�����D$X��� ���  ~�D$���D$������A��� �|$T��   �� �D$�<(��    �$ȍ������D$��T$ �D$X�
   �����0�D$ ��@.�D$fǄ
�   �$ȍ������4�T$��   �L$��ʋD$��  �4$��  ��`  �0   ���4$ǆ�      ǂ     �D$���  �C�T$�r�t$�����1��m�����    �$ȍ�����fǄ(� � �5� �t$�<.�D �F���P��$�  ������PS��E ���   �$��E ���   �t$X�XZ��E ������R�t$\�Pd������������v UWVS��,  �xm  ��m�  ����  �> u��,  [^_]Ð����1���WV��E �Px����t]��WV��E �Px������  ��V�|$,W��E �Pd����W��E ���   ����  �<$��������,  [^_]Ív �������PV��E �Px����u�����W���PV��E �Px�����i����������PV��E �Px�����J����������PV��E �Px�����+����������PV��E �Px������������#���PV��E �Px�������������(���PV��E �Px����������1�|$ ����   �F1�|$ ��$   �t$��5����t$�|$��}�|$�|$�4/��_e����   �J���?��   �ɋ��(������f�����,���P�|$,W��E �Pd�����|$  t@�8 u��F@�P����u��  �R������z{��`t~f���l$���t@���   �c����|$Ƅ,    ��������PW��E �Pd�����|$  t	�v @�8 u���$   ��t���$   A@�P����u��  ��������~t��v �%�   �|$�t$�u�����ɊL �L$�|$��<   �����L ��4   �D����+�7����v VSR�j  ��x  ��������~3H�����������������  P����  V��E �Pd�4$�������X[^ÐVSR�3j  ��(  ����������  J9�~3@�����������������  P����  V��E �Pd�4$������X[^�f�VS����i  ���~  ��E ��F���R����  V�Pd�4$�U�����[^Ív �i  �~  ����������   ���Q��������(/ �	ʉ��������H/ � Ɓ    ǁ�     Ǆ�0     ����  � ���   � ǀ�     ǀ�\     ǀ(�      ��E ��\���Q�������Rd���f�Ív UWVS����h  ���}  �D$0����   9�������   ��(/ �	ʉ���ʍ�(   �M ����0 ��(/ �4 Ɖ��������H/ �>��R�T$��������E �PdZY��7   P���   W��E �Pd��3�0 �E ǃ�     ǃ�\     ǃ(�      ���T$�: u	��[^_]Ð���8 ��`  ���  ��t��R�T$V��E �Pl�����T$t�ƌ  9�uσ�R�~�����묐����   VW��E �Pd��  �     ��(  �  ǃ�     ǃ�\     ǃ(�      ���\����UWVS��(�{g  ��p|  �|$<����  V��E ���   ���G��� w���(�����ᐍG���^��  ��[^_]Ã�V��E ���   ����  ����~ۅ�~׍J�9�~�D�ϊ
�J�B9�u�������  ǃ��      �f���[^_]�P����'���땐��������~���(/ �J�9���  �D- �������H/ ���<���������t����l$�͐���  �c   ����  9�u��l$��������U�[����������v 1�����  ��������  �������V��E ���   ����  ǃ��      �������ǃ��      ǃ��      �����v ����  �������H����  ǃ��      ������(   ���xS��|�����V��E ���   ����  ��9��Y���@����  ǃ��      �C����v ��(   � �2���f��    �%������V��E ���   ��=�   ��������  9�}��.�T$�P��H9�u��T$���.E����  �D ǃ��      ������������j���(/ ����f�VSP��d  ���y  �t$�%�������E V�������Pd�4$�V�����[^�UWVS��<  �d  �y  �D$��$P  ��$T  ����$X  ��   ��<  [^_]Ã�?S��$X  u�F�����  �F؃��  �F�����  ���  ��w����D$��������������랐��$X  u��\$��(   �8����(�  ���v�����H�  �D$��1ۍv �B��D)�9�|B9�|���
9�|B9��  �C��  9�ú�<  [^_]�f��������������)Ћ|$��������<�<���9���9��/  9��Q����L �L��������9�q��~l�k�9�}A� ȉ���ȋt$��H/ ��ډ���򍔑t������  �c   ����  9�u�D$��������(/ 9�|�C��t$��(/ �v ��P�\$��������H����\$�*����:�����    �D$��؍����D�t$��D$� �t$��E �Jh���]  <h�H  </�Q  �D$�x/�D$����  �E ��  ����  ���f�B����F  <:u�r�B����t�ψ��F���t��#��w����t��)���   ~��   PVU��$<  W��Ƅ4@   �D$ ����D$��E �Hh��/�j  Ph�   W�t$<V��Ƅ$?   �,$�D$��E ���   �D���9�r	�'f�H9�t �8/u�9�s��V�D$��E ���   ����V�D$��E ���   ��=�   
�D0/�D1 ��V�D$��E ���   ��X�t$�D$��E ���   ��=�   ���t$�U�D$��E �Pd��Ƅ$/   �|$0/��   Qh�   VW�D$��E �PhƄ$?   ���D$��؍���؋t$��  ���T  ��W�t$����  S��E �Pd�$�������������Ƅ$0   �Jh��$0  Ph�   W�t$<V��Ƅ$?   �4$�����\$���������\$���������Wh�   �D$�������t$<V��Ƅ$?   ����$0  �����|$1u�����|$2r�����|$3l������|$4?������T$5��������L$5�	A��������ЊQ<qu��=u�i�   ��$/  �D$�V��E ����  <&��  ��   ��  �M<%�j  E�L$�1F��f��\$�[����������W�\$�E����������D$�xt��   �D$����  �E �������Ƅ$0   �Jh��$0  �/���Ph�   U��$<  W��Ƅ$?   �D$ �����������u	�B���t<:u���)�x���   ~��   RWU�t$<V���D<@ �4$�l$��E ���   ��Y�t$��E ���   ���=�   PP�t$�W�D$��E �Pd����$0  �Y����xt�����xp����Vh�   �t$�����D$����  �E �������Ƅ$0   ��$0  �/�����������U��������L$-�T$.1�1ҍD$-�D$�\$���D$��XЀ�	w6��0	�u�   �ݺ�   Ƅ0   ������\$��4/  ��F������X���w��W	����X���w���7	�뱐UWVS���K]  ��@r  �D$(��E ������R�������Pd��H   �  ���   �  ǃ0:     ǃ�;     ǃH=     ǃ�>     ǃ`@     ǃ�A     ǃxC     ǃE     ��H/ ��H	  ���v �  ƀ    ǀ�      ǀ�      �  9�u�ǃ�0    ����p���W��H0 P��E �Pd��I ��=  ��  �P��I ������Ѝ��(I UhD  j V��E �P\�    ����I ��������������������hX  h   ��x���P��E �P<�Ń�������P����  V��E �Pdǃ��     XZW�FP��E �PdY_������P�F<P��E �PdXZ������P�FlP��E �PdY_������P���   P��E �PdXZ������P��   P��E �Pdǃ��     Y_������P��  P��E �PdXZ������P��<  P��E �PdY_������P��l  P��E �PdXZ������P��   P��E �Pdǃ��     Y_������P��  P��E �PdXZ������P��<  P��E �PdY_������P��l  P��E �Pd��E j jVU�PX1���,[^_]�f�1��R����VS�t$��t&�D$�T$��f�@B9�t��8�t���)�[^Ð1�[^Ív UWVS���/Z  ��$o  �t$0��tr�L$4��tj���t$<���a ���   ��Z�t$@���a ���   ��)�x=1��ŉ|$��v F�D$9�'�|$0�PU�t$<W�Q�������uމ����[^_]�f�1���[^_]ËD$�L$��u	�f�9�t
@���u�1�ÐS���zY  ��on  �D$���] ��uoǃ�]    ���a ����(���R���h@  j ���������a �P\��H[ �     ��(R �     ǃ�]     ���a �������T$ � ��[����t� ��t�� ����T$��[��f���[Ív VSR��X  �m  ��H[ ���0�����a �t$�ҍ�h[ ��P�Qd����L$$�L� @���X[^�f�UWVS���wX  ��lm  �D$0�D$��H[ ���~N��h[ �D$��1��
f�E��$9.~4���t$W���a �Pl����u��D� �T$�D� ��t��[^_]���v ��[^_]�S����W  ���l  �T$�D$��dt@��etS��x9��] ��[�f������ ����D���] P�1�������[Ð��������P��������[Ð�������P��������[ÐVS�L$�t$�\$1����f��@9�t���u��� [^Ð�� [^�UWVS��@�3W  ,l  �D$�\$Tǀ�]     h   j ���] �|$(W�ǋ��a �P\���; �5  ��������|$$������D$(��] �D$�f��]�} �  ���t$,S�\$�z����Ń�����  ���t$0P���^�������t��p���] ����  �S���] �P����  �����D$�1��f�F@�T����t
��"t��u����߉\$ ؋L$� ���\$��%���PU������D$ �����M  9��4�����-����D$߉l$,�f��D$��8�   ���D$9��  ���t$ V�\$�����ƃ�����   9D$��   �D$��8�   ����   ����3���PV�R���������um���\$��;���PV�5����������p����P���e����D- �(���D$ ËD$�1���v ���?���@�T�T���.�����"u��$����P��t��\- ����D$ ËD$�1��@�T�T���b�����"�Y�����u��O����l$,�]�} �������<[^_]�1��n���U��WVS��L�T  �Úi  �E��(R �M��    �8 ��  ��@����}���^����M���HR �}���E�� �B	�z	 �b  ���u�P���������K  ���u�P����������4  �p����F���PV����������  W��)��~�   �E�RV�}�W�q���Y^��M���R�E�P����������   ���u�P����������   �p����V���PV�j���������   �Eċ ���(����U���W�����M��P���a �Pd���U���)�=�   ~��   �U�PV�Eċ �����M��D P�����XZ��`���PW���a �Pl�����U���������Eċ �����M��D P�������U�������e�[^_]�UWVS����R  ���g  ��(R ���~N1�1ۍ�HR �D$�f�C��   9~1���t$8�D$�P���a �Pl����u׋D$�D ��[^_]Ív 1���[^_]�f�UWVS��   �dR  ��Yg  ��$�   ��m���P���a ��4$���a ��������,$���a �_XV�|$W���a �Pd�<$���a ���   ����~�|�/t����3���R�P���a �Pd�����a �pd��W���   ZY������R�P���$   ���a �P�ƃ�����   Ph   j V���a �P\��h�  VW���a �P ����~>� ��V�����4$���a �P���a �������$����   �Č   [^_]Ð����x���P���a ��<$���a ��,$���a ����a �4$�P��1��Č   [^_]Ã����a ��P���R���1��܍v S����P  �e  �L$���a ��t#��t���] ��~������S���] PQ�RX����[�S�P  �e  �\$�T$�L$���a ��t�@L��t�\$�L$�T$[���[�f�S�UP  Ne  �\$�T$�L$���a ��t�@L��t�\$�L$�T$[���[�f�UWVS��8�P  ��e  ������P���a ����a ������  ��(E �|$Ǉ�      ��h   �P�ƃ����g  Ph   j V���a �P\��j@V�G(P���a �P(������  �D$    ���a �������|$�������|$�t$�T$f��> ��   ���t$V�Pl������   �~0�����a ��u7���t$�L$���   U�Pl�����  ���a �L$���    ��   �L$���  ��?F�i�T$���  ��V�,	����T$���   Q�Pd�T$Չ�$  �F(��(  �����a �D$�T$��@9T$�.����t$��V�P�D$ǀ�   ����ǀ�       ���a �������$�����,[^_]Ív ��V���   �D$,�,$���a ���   ��9D$�y�����U�L$()��P���a �Pl�����W������a ���������a �_����VS����M  ���b  ���a ������R������a h   j ��(E V�P\�    ���a �������$���[^�f�UWVS���M  �ƀb  �D$ �l$$�|$(��(E �   �C    ���a �Rd��tb��P�CP�ҋ��a �@d����tX��U�S(R�Ћ��a �@d����t6��W���   R�ЋD$<���   ƃ�    ���������[^_]Ð������떍������������VSQ��L  ���a  �t$�t$ �t$ �t$�t$�!�����(E �@   ����t���a �t$�   �D$�BdZ[^��f�X[^�UWVS���L  ��la  ��3���S��(E �n(U���a �Pl����t=��U���a ���   ����~-�P��|'/u�E�Ht)�T(��/u��D( ���������[^_]�u�V)�����u���S�F(P���a �Pd����f��D' ��1�븐WVS��K  ���`  ����(E �~(W���a ���   ����~ �|'/t����3���R�P���a �Pd�����a �xd����(V���   ZY�t$�V���D�����[^_ÐUWVS��   �TK  ��E`  ��(E ���   ��x;��  �  ���C(P�l$U���a �Pd�,$���a ���   �ǃ����  �|/t6����3���R�T$U���a �Pl����t���T$R�W���a �Pd���{��tb�����   W���a ���   ����t7���a �pd��U���   ZYW�P�֋��   ����t	��U�Ѓ��    �Ĝ   [^_]Ív ���   ��x�;��  }����a �pd��U���   ��XY�?������   P�R�f�� �����$  ������������   P���������f��!�������3���PU���a �Pd���{�������c����v UWVS��,�I  �à^  �|$@�t$D��(E �E ���C  ���a ���[  �L$H��p������T$����L$�T$L���������1�T$��jh   @h,  h�  �LQ�L$ �TR�PT��jh����h,  h�  �t$,V�|$$W���a �RT��h����jh�  VW���a �R@��h����jh�  ��,  RW���a �R@��h����h,  jVW���a �R@��h����h,  jV���  R���a �R@�|$(��
��jh����jj�V
RW���a �RT�t$4���� h   ������RV�D$�PR���a �RDh   ��URV�D$$�P2R���a �RD��h�   hfff��U(RV�D$$���   R���a �RH�t$4��(�� �}��  �D$
   ��   ��j�P�D$h|  VW���a �R@��h����jh|  VW���a �R@��h����jh|  �D$�PW���a �R@�D$4��*�� 1�������L$������L$�|$���g�v �L$�D$��jjW�D$�PRQj ������ h   ��D$������   P�GP�D$��#P���a �PD�D$�D$�����L$9�td�t$��   9��  ~R9��   u'��h�׳�jhz  �G�P�D$$��P���a �P@�� �6�0����$  ���C����L$�>���f��D$��  �}��   �L$�D$���   h   ������RW�t$�VR���a �RD�D$$�   �t$��<�$����jh�   P�D$ V���a �R@��h   �jh�   �D$PV���a �R@�� h   ����   RW�t$�VAR���a �RD���L$��jh����jj<Q�L$ �|$$���   R���a �RT�t$4��  �� h   ������RV��  R���a �RDXZjh�z �jj<�L$Q��@  R���a �RT���a �RD�� �}t<������j�PV�D$O  P�҃��   ��,[^_]�f��D$   ��   �G���f���������1���,[^_]�f��"E  ��Z  ��(E � ��t1����a ����Ív UWVS����D  ���Y  �T$8��(E ���tg�D$0-�  ��9�S���  9�|I�|$4��,  ��;|$<7��,  ;t$<|+�p	9���   �p(9�|)�w	;t$<} �w;t$<|�����f��   ��[^_]Ív �q�t$N�
  ��   ��|  9�|�o(9l$<|v�;t$<|n�T$<)�����������   x�9��  ~�9��   ��   ���   �|$u�k�0��$   �x���PP���a ���   R���   R�Pd���V���f���  ���   9�},��6  9�|"9t$<�0�����  ;l$<|�    �������?  9��
���|  9������9t$<�������  ;|$<������������������   �����k�0��$   u�|$ �>����у����   P�4���������S���C  ���W  ��(E ���t�|$tn�|$
t�{t�   ��[Ív ���e�����v �����a ���   R���   ���|$t0�L$�Q���^w���>��L$���   Ƅ�    �f��    뗅�~�Ƅ�    �f�S���u�/�v 8�u@�Z���t�ڊ��u�1�8���[Ð�Z1�8���[Ê��VS� B  ��W  ��� ���   S�A��� ����ȍ��� ����  �  �@ ��9�u����ȍ�ǀ�     ǀ�    ��[^Ív ǀ�    ��� �u�O�������ˊH@B�Z���u�� 1���[^�UWVS��P  �tA  ��eV  �t$�D$�B�$�B�r�t$�v 9$~3�*�t �t$��� t
�s����wp@�B�\$�;
tK�B9$Ѝv �D$��$H  �B��$L  �D$@    �D$D �t$@�D   �|$�D$��P  [^_]��D$�\$�Z�B   �q������t���/�u  �p94$�i  �|5 ���/��   ��*�Q  �r�\$�;
�
  �r�N�J�p�r�?
�  A�J94$��   �\��v 9$�/����;/��   C�ƍF�B�K���
tu�z�o�j���������*t�9$u���������r�|5�
t3�z�O�J94$������D5 <
��  ����  F���r�|5�
u��D$�\$�Z�   ���v �D$�|$�z�B   9$�_����H������A�����F�B�;
�Y  ���z�&���f��D$�t$�r�   �J�p�r�?
������D$�L$�J�   ������D$�t$��$H  �Z��$L  �| ��D$�������D$�HЀ�	��  �D$<"�U  <'�M  �D$����߃�A����   �D$@   �$A�ϋD$)ǻ   �t$C�4$9�t6�t ���߃�A���  ���_�  ��$�  �NЀ�	��   �DC �D$�������v��&����|$D����u��   �8�u@A�����   ���u���F�����   ��̋B������D$�t$�r�B   �����<_�0����|$$�%����   �D$<�D$�T$ ��݉ËD$ȋ4$9���  Iu�T$ �D$@   �D$@�B�<
��  �M�J�D$D�D$E �t$@�D   �|$�D$��P  [^_]�@�B�L���
��   �rF�r�4$�C�����9 �����D$@   ��D$@   �$�t$)�1�1ۍL$C�L$�L$�$���iЉ�<	�D  �4���t�C�D$��J�L���
tD�B�h�j�D$��$9�u��$�DD ��$D  �t$@�D   �|$�D$��P  [^_]��B�   ��B�   �.����t$F�r��D$<
t{�C�B�D$@   94$��  1��D$C�D$�l$�D$�0�8D$��  ����  �N�J�<
tA�Z�k�j<\u>9$�_  �D$Ȁ8 ��  G�D<C\��몋D$@�B�   �v����B�B   G�t$�>9$��D<D �;����D$<    �T$1��t$�@9�t��@9�u��D$<�D$�D$�������+��N����|$,�L$$�\$(�\$��t*�ً|$�f�8�uG@����t��u���F���tl��҄�u�|$$�T$ �l$(�D$@   �D$�L$D��t�\$CA�A����u�� 1ɋD$�4$9�}�X�Z�| 
t)�BA9��b����B�4$9�|���|$,�L$$�\$(�����B�B   ���D$D �/����������G�D<C\������L$A�J�   ������l$�D<D 94$������F�B�|5 
tJ�B������N�J� <
tS���Z<rtB<tt7<n�p����
�i�����l$�D<D �|$ t������v �B�B   �����	�:�����3����B�B   �
�"���f�WV��  �ǋ�4  ��t�G��  ^_É�����m����G�D   ����  ^_�WVS��  �Ë�4  ��t'�{��$  �D   �ǃ4      ��  [^_Ív ��ډ������{�D   ��  [^_Ð�D$�O�����t�     ËD$�;�����t�    ËD$�'�����t�    1ҋL$���P�f��D$������t�    �T$�PÐS�\$�D$�������t �    �P���t�v CB�J����u�� [�UWVS��<  ��8  ���M  �D$�ӉL$��t	�:��   �D$    ��$P  ��t��$P  �8tu�D$    �D$�����  �ȋl$��N����+�8���   EG�E ���t��u�8���   ��t�;t@���D$ �\$�P�t$�����������<  [^_]Ð�@�D$늍v �B�D$�\����S�K�|$0����tB@�H��
��u��  ��$P  ��t��$P  � ���%  ���7  ��W�t$����������<  [^_]Ív �ʋl$��Q����-f�8�uEG�U �����   ��u�ʋl$�*��������8�uEG�U ���t��u�8�tw�ȋl$��3����/�v 8�uEG�E ���t��u�8�ub�\$��t�D$����D$���t$�t$�����������<  [^_]�f����s������D$ �\$)��������D$ �\$�������ȋl$��*����%�8�uEG�E ���t��u�8�ud�\$��t��D$����T$�s�����$P  �@�D$/ ���
  �D$.0�0�   �T, ���|$0 t	�@�8 u�f�B@�H��
��u��  �}����ȋl$��4����=�v 8��6  EG�E ���t��u�8��  ����  ��$P  ����  ���$P  ;��   ��t����  ����   ����$X  �@9C����P�t$���\������|�����$P  �H���|$0 t�@�8 u���$P  �S���3���A@�P����u��#�����y�ۺ   �L$!�L$�D$�|$�׍v �|$O�ع
   ����J0���D$�8����������u׋D$�|$����   �l$������j �t$��������������ʋl$��,����=8�uEG�U ���t��u�8�������ʋ|$��0����!8�uGE��E ��t��u�8���   ����   ��$P  ����   ���$P  ;��   ��t����  ��u}PP��$X  �@9C�������D, -�-�������;�$X  ���q�����$P  �H�{�C��$P  �S��u�8�uG�Q���t�ъ��u��8����.����Q���j�t$������������QQ;�$X  ��� ����|$��3����!8�uG@����t��u�8������������D$�*�������  ��^����D$�������r  ��7����D$��������I  ��:����D$������Ņ��  ��=����D$������ǅ�tt���������t	�������{ �������$P   t&��$P  � ��t.��u��$P  �x ������RRU�t$���r�����������$P  �h�ލ�@����D$�C�����tl��t���t��u
�{ �������$P   t&��$P  � ��t.��u��$P  �x ������PPW�t$���������������$P  �x�ރ��t$�������������QQ�\$9\$ ���L���SS�\$9\$ ���:���WW�\$9\$ ���(���UU�\$9\$ ��������$P  �P�C�c���RR����������v S�1  �âF  �D$�{�����tB�    ��� ��?1�H��� ������ȍ��� �B��H  �  �@ ��9�u��[Ív S�I1  ��>F  �D$������t?�    ��� ��?.�H��� ����ȍ���a �B���   �  �@ ��9�u��[�f��D$��t��  Ð�D$��t��  �Q���  ��~��     ÐUWVS��<�0  �äE  �t$T��t�>w����H���������N���P�t$\�i�������<[^_]�f�����]���P�t$\�I�������<[^_]�f�����X���P�t$\�)�������<[^_]�f��F��tm��C�����P�t$\��������<[^_]Ív �F�D$/ ��uH�D$.0�   ���D,P�t$\���������<[^_]�f���V�����������<[^_]�f���H���둉�x\�   �|$�D$�|$�v �t$N���ȿ
   �����0�D$�0����������u׋D$��x�l$�p���f��D4-�d���f����UWVS���C/  ��8D  �t$$��t���tG��tZ��t��j �t$,���������[^_]Ã�1��V����P�t$,���������[^_]�f���V�����������[^_]�f��V�F< u	f�B�< t�<-tI�
�A�1�<	wV1�D� �4 �A����,0B�
�qЉ�<	v��t�݃�U�t$,�M�������[^_]�f��r�J�A�<	w��   �f�1���VSS�K.  ��@C  �t$��t���tww!��t\��t7��j �t$�������Z[^�f�����w��j�t$������Z[^Ív ���N������P�t$������Z[^Ð��V���������Z[^�f����~ �ˍv UWVS���D$ ����   �8��   �@����   ��@  ����   �Ƌ|$$��\$1��$f����T$$��u�   �v 8�uC�J���tb�ʊ
��u�G��D9�u΋$��@�������T$��t�\$$CA�Q����u�� ��@  ����ы|$(�|�@B��@  ��[^_]�f��B��u��$������|$(�|�@��[^_]ÊD$�܋|$$��\$냐UWVS���,  �A  �D$�D$4��tM�8uH�@��tA��@  ��~7��1��D$����T$8��u�\f�8�uC�J���t.�ʊ
��u�G��D9�u҃��t$<�\$��������[^_]Ív �B��uӋD$������D�@��[^_]Ê��f��D$��t'�8u"�@��t���   ���J���   �L$���S����+  ���@  �D$��t �8u�@��t�T$��x�T$9��   ���t$��������[Ð�����v �D$��t�8u�@��t���   Ð1�Ð�D$��$� �  �@ ��9�u�Ív WVS�\$�D$��N ��l�V��N �<�    �7������$ ���t@B�J����u�� ������ǃH$     ǃL%     ǃP%    �D$��T% 1�[^_ø�������v UWVS�t$��$ ��~8��  1�f����tA�L$���f�8�uC�Q���t�ъ��u�G��H9�u�1�[^_]Ív �A��u�F@[^_]ËD$� ��UWVSR�D$��$ ����   ��  �|$��\$1��D$�v ���T$��u�   �v 8�uC�J���tn�ʊ
��u�G��H9�u΋D$��n�T� ���  �T$��t�\$f�CA�Q����u�� ��$ �ҍȋ|$ ��D  ǁH      B��$ X[^_]Ð�B��u��D$���|$ ���D  X[^_]ÊD$�ދ|$��\$�w����D$� �f��D$ǀ�     ƀ�  �f�S���.)  ��#>  j ������[ÐS���)  ��>  �t$�t$�������[Ív S����(  ���=  �t$�t$������[Ív S����(  �ÿ=  j �V�����[ÐS���(  �ã=  j �:�����[ÐS���(  �Ç=  j �6�����[ÐS���v(  ��k=  j �������[ÐUWVS���  �\(  ��I=  �<$�ŋ�4  ����  �@�D$�E���q  ����  ����  �D$� ��tT���Z  ���O  ��$  �D   �|$�ǅ4      ����8  �\$�R����D$ ���D$���  [^_]ËD$�H�L$�P��$p  �D$��t�v A@�P����u��  ����  ��$  �D   �|$�ǅ4      �D$ �D$��t$��������D   �|$�E���
  �v ��8  ��$ ��~R��  1��D$�l$��f������  ��L$�f�8�uC�Q����.  �ъ��u�G��H9�uʋD$�l$��N ��~]��$ ��$p  �\$1��D$�l$�͍v ����6  ��T$�f�8�uC�J�����   �ʊ
��u�G��P  9�uǋD$��P�\$������D$ ������f��t$ �t$��������}�D   �E�D$�E����
  ��4  �����������  ��t$�������D   �|$��  �t$ �t$����a����D   �|$󥋅4  ��������d����v �A��������F@�D$�D$���  [^_]ÊB�������D$�l$��P�\$�����ǉD$ �    +�8  �����������ʉ���)��ȍ�������؉G���t����E�D$�}���������t$�$��C����t�v 8��}  FA����t��u�8��g  ���  ��$  �D   �|$�ǅ4      ��j��8  �\$�k����D$ ���D$���  [^_]ËD$�x�|$�x����������t$�(�$��v����8���  FA����t��u�8���  ����  ��$  �D   �|$�ǅ4      ���T  �D$��4  ����  �}�U����D$�P���F����$��~����)�\$����-���8��%���CA����u��������4  ����  ��$  �D   �|$�ǅ4      ������t$ ��������D   �|$��������t$�$��H����ff�8�uFA����t��u�8���  ���t$�n�$��X����8�uFA����t��u�8��  ���t$�$��N����u�8�uFA����t��u�8������t$���$��&����v8��:  FA����t��u�8��$  ���5
  ��$  �D   �|$�ǅ4      �D$ �D$��t$���#����D   �|$󥋝4  �E�}��  �Ǆ��d����t$�i�$��s����8�uFA�����8
  ��u���t$�w�$��x����T$�߈��8�uF�D$�D$�� ���  ��u���r�<$�������t$�������8������FB����u�����������  ��$  �D   �|$�ǅ4      ����  [^_]��  ��t$���[�$�������v 8�uFA����t��u�8��  ���t$�{�$�������8�uFA����t��u�8��  �t$���!�$�������8�uFA����t��u�8���  �-�4$��Q����t$���������8�����FB����u�����������  ��$  �D   �|$�ǅ4      ���k�����t	�8��  1���P�&f���$  �D   �|$�ǅ4      ����  ��8  �\$�U����D$ ���D$���  [^_]Í�$  �D   �|$�ǅ4      ���EP��8  �\$�*����D$ ���D$���  [^_]Ê�$p  �_�������  ��$  �D   �|$�ǅ4      ����8  �\$�����D$ ����������  ��$  �D   �|$�ǅ4      ����8  �\$������D$ ��4  �ǃ����4  �U�$�������D$��$p  �D$������
  �D$�@��t �t$�}�L$8�uFA������  ��u�|$�|$�   1���tj�U����  �   1��|$����wۋD$�@����  �L$�T$�AB�B����u�� ���"  ��$  �D   �|$�ǅ4      �t$ �t$����.����D   �|$󥋝4  �U����  ���l�����t$��������D   �|$󥋝4  �U���B����E��������t$�,�<$��������������8������FA����u����������J  ��$  �D   �|$�ǅ4      �D$ �D$��t$���j����D   �|$�U��4  �_����t$ ����D����D   �|$�������t$ ����'����D   �|$��X����D$�@���������|$�4$��
����:�v 8�uGF�����-  ��u�������D$ �D$��������������m����t$ ��������D   �|$��U����|$�_�\$����  �L$�t$�<$��v����|$���(8�uFC�����.  ��u�\$f���������C��������t$�.�<$��������v ���l���8��d���FA����u���R�����4  ����   ��$  �D   ���ǅ4      ��t$��������D   ���E���m����D$��$p   t	�v @�8 u�f� . �D$��$p   t	�v @�8 u��S��t�L$�v A@�P����u��  ��4  ��td��$  �D   ���ǅ4      ��t$���B����D   ���E��������t$���#����D   ��󥋅4  ���?����$����v ��t$��������D   ��󥋅4  ��u��f���4  ���������t$��������D   �|$����������������  ��$  �D   �|$�ǅ4      ���  P�t$�t$��8  �\$�7�����4  �����o��������D$�@���>������U����0�����t$ ����+����D   �|$󥋝4  �h������  ��$  �D   �|$�ǅ4      ��j ��������  ��$  �D   �|$�ǅ4      ����8  �\$������D$ ����4  ���-  �E�<$�������|$�|$ �|$��u1�D$�@��t&�\$�]�L$8�uCA����t��u�8������f�����  VP�t$��8  �\$��������4  ����   �}u͋D$�@����t��t$�<$�������,��v ���z���8��r���FC����u���`�����4  ��tZ��$  �D   �|$�ǅ4      �\$ ��������D   �|$���E������t$�������D   �|$��S����\$ ����i����D   �|$��󥋍4  ��u�럍t$ �t$����?����D   �|$󥋝4  ��������U�,����t$ �t$��������D   �|$󥋝4  ������������v �D$������t$ ���������D   �|$�� ����T$�X����t$ ��������D   �|$���������������i  ��$  �D   �|$�ǅ4      �D$ �D$��t$���`����D   �|$��}�}�  ��4  �����c�������f����������4  ����  �L$�(�T$�\$�������8������AB����u���������4  ����  ��$  �D   �|$�ǅ4      ��t$�������D   �|$�1��1�C���8  ���,  ��4  ����   �}��   ����  �D$�8u��x����t��t$�)�$��~������t�8�u�FA����u��u������b  �)�<$��~����t$8�uFB��
��t��u�8�9  ��4   ��	  ��$  �D   �|$�1���4  �  ��t$��������D   �|$��8����D$�P���3����t$�$�������,�������8�����FA����u��� �����4  ���g  ��$  �D   �|$�ǅ4      ��t$���G����D   �|$������t$���l�$��E���8�uFA����t��u�8���������t$�c�$��m���8�uFB�����  ��u�����������  ��$  �D   �|$�ǅ4      ���������t�����  ����  �   ��P�@����t$ ��������D   �|$������t$ ����d����D   �|$������t$ ����G����D   �|$��r�����$p  �D$�����t$ �t$��������D   �|$󥋍4  ������������t$ ���������D   �|$��b����t$ ���������D   �|$󥋽4  �����t$ ��������D   �|$��c��������������t]��$  �D   �|$�ǅ4      �D$ �D$��t$���]����D   �|$�M�}��  ��4  �����������f��t$ �t$��������D   �|$󥋕4  ��u�랍t$ ���������D   �|$��0����@�������D����D$�8�y  ��$p  ����  �ʰc�   8���  �D$�0F�$�������t��u�8���  ����$8  PS�\$�����D$ ���$�������  �L$��$p  �|$��AB�B����u�� ����   ��$  �D   �|$�ǅ4      ����8  �\$�����D$ ����4  ��tu�}�B  ��8  ��$ ��������H��$ �4�    ����  ��$p  ��t�|$GC�K����u�� ��ʋ|$��D  ǀH      �B�����t$���|����D   �|$��n�����t$���_����D   �|$��.�����t$���B����D   �|$󥋽4  ��������c�����t$�������D   �|$�E�D$������������������ʰc�   8�u�D$�0F�$�������t��u�8��6����Ⱦc   �<$�������|$�L$��8�uGB��2��t���u�L$8��  �ȋ<$�������c   �|$�L$��8�uGB��2��t���u�L$8��  �ʋ$�������|$�8�uGF���t���u�8��  �ʋ$�������|$�8�uGF���t���u�8��  �ʋ$�������|$�8�uGF���t���u�8t+�ʋ$�������|$�8�uGF���t���u�8�Z  UU��$8  PS�\$�����D$ ���=�������  �ȋt$�(�<$��v���8�uFB����t��u�8��  ��4  ����������  �\$�(�4$��v���8�uCB��
��t��u�8��   ��4  �4�����t$��������D   �|$󥋕4  ���e�����������y������������t$ ��������D   �|$��Y����t$ ��������D   �|$��L������3������   �Ɖ�������8��   ����8  �\$�d����D$ ����t����B  ���9  ���*
  1ۉ������8��������<$�������7��������������������  ���  [^_]��	  ���<$��~�����������d������w����X���PP��$8  PS�\$�����D$ ���c���PP��$8  PS�\$�����D$ ���C���PP��$8  PS�\$�"����D$ ���#���PP��$8  PS�\$�����D$ �������$�������t$�8�uFB���t���u�8
��   ��t��$0  �8t2VVj ������~ ���������  �D$�   ������  ������1��k�
�T
�@��YЀ�	v�WWR������@���r����E��������<$��1����=�\$8�uCB��
��t��u�8��������������  �D$�s�����$p  �D$�������x������t$���?����D   �|$��a����$�������L$����&  8��  AF����u���  ��8  ���[  SS��$8  P�\$�����D$ ���������r����E�D$����8  �\$�����D$ ���D$�  �>�}tl���K������t	���;����C���0������`  �D$�L$�����D$�E����  �Ë�4  ��u���t$���;����D   �|$�뎊E��t��t$�<$��~����)8�uFB��
��t��u�8�d����������X����$�������L$�
��ti8�ueAF����u��uW��8  ����   RR��$8  P�\$������D$ ���Y�����4  �����QQ�\$������RP������D$ ���/����4$������D$�����ǋ�8  ��t;��tWW��$8  P���o����D$ �������SSj P�\$�U����D$ ���������N ��$ ��9�������1ۉD$���tRC�D$8D$uG��D$�D$��D$�|$ u؋D$��P  �|$ t*G�UUj P�\$�����D$ ���`����D$��P  G닉�H   �������L  �������QQ��$8  PS�҉D$ ������UWVS��,  ��	  ���  �Ő���a����D$��4  ����  �}�|  �E�D$f��D$�D$�u�����]  �|$��1����=f�8�uGA����t��u�8��N  ��|$�+��%���8�uGA�����&  ��u��|$�-��(����f�8�uGA����t��u�8���   ���|$��+����*8�uGA����t��u�8���   ���|$�/��.���8�uGA����t��u�8���   ���|$�+��N���8���   GA����t��u�8���   ��4  ����  �}�|$��$  �D   �ǅ4      ���������P�L$�T$��8  �l����D$����4  ���  �}������D$��,  [^_]�f����������4  ���B  �}��$  �D   �ǅ4      �����v ���|$��Q����-f�8�uGA����t��u�8��$������|$�*������8�uGA����t��u�8���������|$��3����/8�uGA����t��u�8�������|$����*����%8�uGA����t��u�8���������|$��4����=8�uGA����t��u�8���������|$�=��,���8�uGA����t��u�8��\������|$�!��0���8�uGA����t��u�8��4�����|$��3����!8�uGA����t��u�8�������|$�������<8�uGA����t��u�8���������|$��^����>8�uGA����t��u�8���������|$��7����<8�uGA����t��u�8���������|$��:����>8�uGA����t��u�8��l�����|$��=����&8�uGA����t��u�8��D�����|$��@����|8�uGA����t��u�8�������1����?��t$8�uF@����t��u�8�]����������������Ɖ��[����8�=�������
�����������'������u������b����\$��t�����   ����   �D$�������t$��������D   �|$�������v �t$����s����}�|$�D   ��v����t$����S����}�D   ������t$����7����}�D   �������\$�S�t$���h����f���UWVS��,  �  ��u  �ŋ�4  ����  �}t1���z����$��4  ����  �}��  �$��,  [^_]Ð�E�D$�E��t��t$�������{���t�8�u�FA����u��u���4  ����  �}�|$��$  �D   �ǅ4      ����8  �L����D$����4  ����  �������D$��E��t<���U����������$��4  ��u܍t$���������D   �|$�E��u��u����t\$�}�L$�f���t�8�u�CA����u��u�����������}�L$�\$��������8������CA����u���������4  ���  ��$  �D   �|$�ǅ4      �����t$����C����}�D   ��I����t$����'����}�D   �}�P����M�E���B�����3����;��v ���-���8��%���AC����u��������4  ��t?�}��$  �D   �ǅ4      ������t$��������}�|$�D   ��7����t$��������}�D   ������t$����d����D   �|$��!����t$����G����D   �|$��t����v UWVS��l  �  �Ù  ��$�  ��$�  ��$X  Ǆ$\      Ƅ$`   ��$   Ǆ$$      1��: t	f�@�< u���$(  Ǆ$,     Ǆ$0     Ǆ$T      ��U�����Ã��D$�D$��$   �D$�"f���$4  ��tH�D$�d����Ë�� ��u3��$T  ��uՋT$�t$���N�����$4  �D   󥋄$4  ��u��؁�l  [^_]�S���   �Ó  j j �`�����[Ív S���~   ��s  j j �@�����[Ív VS���]   ��R  �t$V������P��5���PV������4$������P��=���PV������4$�h�����P��F���PV������[^Ë$Ë$Ë4$Ë<$Ë,$Ë$�         \��x��\��x��\�� �����h!��\�� !��4$��h ��X��|���#��0#�����0��h��h��@�����t�������\��\������d����\����\�����������������������t��������������l�����"��0��0��0���!���!��<"��j���i��di��Hi��0j��i���i��i�� i��v���0���0���0���0���0���0���0���0���0���0���0���0���������0���������������������������������0���0���0���0���0���0���0���������������������������������������������������������������������������������0���0���0���0������؃��ă��(���ă��ă��ă��ă��ă��ă��ă��ă��ă��4���ă��ă��<���ă������ă��ă��ă��ă��ă��ă��ă��ă��ă��؄�� ������@���T�������                               �����   �                                                                                         ����                       �                                                              �����   �                                                                                      ����                       �                                                           |�������ܺ�����8�����������rgb black white red cyan magenta silver maroon olive lime aqua teal navy fuchsia purple orange pink brown coral crimson gold indigo khaki lavender lightblue lightgray lightgrey lightgreen lightyellow salmon skyblue tomato violet transparent none solid dashed dotted double groove ridge inset outset html title div span br hr h1 h2 h3 h4 h5 h6 img ul ol li table tr td thead tbody form input button textarea strong code pre blockquote script meta link header footer nav main section article aside figure figcaption details summary label select option < H Search Google or enter URL R background-color background font-size font-weight bold 700 font-style italic text-decoration underline display flex inline-block margin-top auto margin-bottom margin-left margin-right margin padding-top padding-bottom padding-left padding-right padding border-radius border-width border-style border-color border border-top border-right border-bottom border-left line-height text-align center justify overflow visible hidden scroll visibility collapse position static relative absolute fixed sticky z-index flex-direction row-reverse column column-reverse justify-content flex-start flex-end space-between space-around space-evenly align-items stretch baseline align-self flex-wrap nowrap wrap-reverse flex-grow flex-shrink flex-basis gap min-width max-width box-shadow href src alt class target _blank type document.write [ input ] [Button] Untitled Error Loading... www. .org .net .edu .gov .io https:// 0123456789ABCDEF http://www.google.com Enter URL or search New Tab Web Browser File New Window Open URL... Close Tab Edit Copy Paste Select All View Reload View Source Full Screen [FW] cm_init: Done.
 fs_new_folder fs_new_file <Menu name=" </Menu> <Item label=" id=" <key> </key> <string> </string> CamelMenuDef [FW] Loading config for:  Info.clist [FW] Picker Refresh...
 [FW] Picker Refresh Done.
 * [FW] Dialog Init...
 [FW] Dialog Init Done.
 Open /home Save ^ Name: Cancel Out of value slots var % === != !== <= >= && || true false undefined null [object Object] const if ( while ) return , console.error console.warn document.getElementById document.querySelector window.alert parseInt String Number [ { } ! else console.log console.info Boolean += -= *= /= ? ; console document window ++ -- function for do switch case break continue default this new  ________________________________________    Error: Failed to load page

URL: %s http://www.google.com/search?q= [FW] WARNING: cm_init called twice!
    [FW] cm_init: Setting up framework...
  [FW] Failed to allocate config buffer
  [FW] Config not found (or empty):   [FW] Config loaded successfully.
   C   S   G              H       B   ,       9       +   -          7       %      !                            J                Q       A               1           <          L          F      ?   R   :   =         $         '   4   M   0          D                       "      @   I                                *                  .   C                         N       6       ;               
   	   3                       O       K                   >           )                   &                       E              8   #                   (       /   5       2   P   C         	   �� �H*�`
a  JpR���I  �{.�U  )�b   ) ���&                               	   
                                                                   !   "   #   $   %       &   (   *   ,   .   0   1   2   5   6   8   9   :   ;   <       =   >       @   B   C       D   E   G   I   K   M   O   P   A�ze��L�q,��A�\DI�%�Pr���=�ijі+R�j�������p����bϐ��	97(2�� �D���T]�Ѝ���`I��RӭI��P�YD�H.�C��،a5���
�G���@�>�!wp��	�K�d�K/q|M-(��^4iB���Bd8��KJ�H�|���nx�c%1rMw9�!���@M�xy�@�����)X={?7�B�	K��"��h#���ۏigsc�ۗs�>c*�|�c�磦�>Rn7�~�!����� E��(�2�?uz5�^J��	%S�>f��^�Vm+�]�Z�Ӊ;����*`(���$6~��f�    ����                           ��  ��  ]�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  "�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  6�  �  ��  �  �  ��  ��  ��  ��                          ��  ��  �  ��  �  �  ��  ��  �  ��  ��  �  �  �  �  ��  ��  ��  ��  �  #�      @� �r  p   H 4!  ��  �  ��  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   X�  ���o��     \�    ,� 
   �           ��    �              ���o?                                                           ^   �       /  (�  8     C  $�       @   ��  ��    �  D�  :     �  T�  ^     �  �  k     d  ��  v     �   �r  W    �  P�  "     �   �>      )    �  �     �    H @    z  �>  	    `  ��  �    �  ��  V     W   m  O     �  T�       �  (�         T�  �     �  ��  3    C  ��  0        ��  @          |     �  <�       �  t�       M   DX  �    n  @�       �  ��  !     �   Lz  �    �  �  a       ȋ  {     �   p  �    �  H�  
     �   �G      u   �n  s    v  \�  �     �  �1      �   0}  5     T  ��  �    r  0�  �    [  ��          4!  H    �  �  l      �  �     p  ��  �     �  Ю       �  l�          �  �     �  ��  4     �  �  :        ��       Q  ̫  Q       P�  �     �  Ć  D     I  ��  %     �   h}  �     �   �~  N     �    ~       5  �  �     8  �  �    &  �       '  �  �     �  Ċ  \     �  T�  �     S  ��      l   �m  5     �  Ħ  #     <  `�  �    �  �  �     4   ��       �   �r  8     `   hm  V     �  ��       '  D�  �    �  ��  !     
   @�      p  �         �       �    ~  �     �   �m  �     �  <�  c      on_paint current_url status page_offset page_title content_len page_content fetch_url nav_back nav_forward nav_home switch_tab on_input open_url_new_tab on_mouse cdl_main my_memcmp my_strstr my_strchr cm_init actions action_count config_count cm_bind_action execute_action_by_id internal_menu_callback strncpy_safe parse_menus_from_string parse_plist_xml cm_get_config cm_load_app_config cm_apply_menus cm_draw_image cm_draw_image_clipped cm_picker_refresh cm_picker cm_dialog_init cm_dialog_open cm_dialog_save cm_dialog_up_dir cm_dialog_select_dir cm_dialog_submit cm_dialog_render cm_dialog_handle_mouse cm_dialog_click cm_dialog_input js_new_undefined js_new_null js_new_boolean js_new_number js_new_string js_new_object js_new_array js_value_ref js_value_unref js_to_string js_to_number js_to_boolean js_object_set js_object_get js_array_push js_array_get js_array_length js_init js_register_native js_get_global js_set_global js_get_error js_clear_error js_console_log js_console_error js_console_warn js_document_getElementById js_document_querySelector js_document_querySelectorAll js_window_alert js_eval js_window_setTimeout js_window_setInterval js_register_dom_api   ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��      �     �      �     $�     (�     ,�     0�     4�     8�     <�     @�     D�     H�     L�     P�     T�     X�     \�     `�     d�     h�     l�     p�     x�     |�     ��     ��     ��     ��     ��     ��     �d       D|	  4           /}      %�  %�  �  -   R  L   Eq	  	Z   
_   y   y   y   y   y    Fint !  
�   
�   �   y    �  �   
�   �   y   y   y    h  �   
�   �   y   y    *0  �     I  ##       -    %�  G    3  -    2 d  �  
d   �  4t  �  	y   �   t  -    �   �  -    �  3  *�	K  �  [   F  v    �  �  �    �  1   �  �  !�  E  "�  �  %
   �  &
  $�  '(  (�  (A  ,r  )�  07   *�  4�  +�  87  .n  <-  /�  @�  0�  D�  1�  Hn  2�  L�  3  P[  4<  Tz  5`  X@  8z  \�  9�  `�  :�  d�  ;�  h*  <�  l�   =�  p�  >   t   ?  x*  @�  |7  A3  �Y  BG  ��  C\  ��  Ff  ��   Gf  �  Hf  ��  I�  ��  Jf  �  M
  �E  N�  �h  O�  �  P�  �  Q�  ��  R  ��  S>  �K  Ta  �1   Uu  ��  V�  ��  W
  �   X
  ��  [�  � V  V   
  
K  L   o  o   %�  
`  L   �  L   o   
{  �  L    
�  H
�  y   �  V   
�  y   �  V  V   
�  �  �  y    
  
�  y   
  V  �  y    
�  y   (  V  L   y    
  y   A  V  y    
-  @   n  V  y   y   N   �   �    
F  �  y   y   y   y   y    
s  �  y   y   V  y    
�  �  y   y   V  y   y    
�  �  y   y   V   
�    y   y   y   y   V   
�  <  y   y   y   y   y   y    
  [  @   [  y   �    
�  
A  z  L   y   o   
e  �  L   �  o   
�  I
  �  �  V   
�  �  �  V  o   
�  y   �  V  V  o   
�  �     V  y    
�  �    V  V   
  y   3  �  V  J 
  o  G  V   
8  \  y   �   
L  K4   
a  �  �  �  �   
y   
k  y   �  y   y   y    
�  y   �  y   �  y    
�  y   �  y   �  o  y   �  y    
�  y     y   �  o  y    
�  y   >  y   L   o  y   L   �   
  y   a  y   L   o  y    
C  y   u  y    
f  y   �  �  �  �   
z    ]�  *$_	�  �  _#   "  _'L     �  _3�  *,`		  �  `#   �   `)y    �  `6y   $�  `R	  ( 
�  :	  `]�  
	  
�  %�  %�  %�  %�  %�  %�  Lsys (	  �1   y	  -   ? *�C	�  �  D4    �  E4     F	y   �  G	y   �  H	y   �  I	y   �  J	y   +  K	y   E  L	y    U  M	y   $  N	y   (�  O	y   ,:  P	y   0q  Q	y   4�  R	y   8�  S	y   <�  T	y   @T  U	y   D|  V	y   H,  X	y   LE  Y	y   P  Z	y   Tx  [	y   X�   \	y   \)  ]	y   `  ^	y   d�  _	y   h'gap `	y   l�  a	y   p  b	y   t  c	y   x�  d	y   |�  f4   ��  g	y   ��  h	y   �  i	y   ��  j	y   �t   k	y   ��  l	y   �  m	y   �b  n	y   �   o	y   ��  p	y   �H  q	y   �x  r	y   ��  s	y   ��  t	y   ��  u4   �   vy	  ;-   |!  v   @  '  �   �  ��  ;-   ��     
  �  x  �  [  H  B  S  \  	�  
�  �  �      �  d  �  �  �  
  c    �  #  �  �  �      0  1  �   p  !!  "�  #�  $  %d  &:  '�  (L  )�  *�  +�  ,�  -R  .�   /�  0�  1�  22  3k  4f  5   6�  7�  8 7  �-  M�  D��  A  �!   <  ��  �   �
#  �  ��  (R  �	y   ,=  �
�  0)src �
�  0)alt �
�  0)id �
i	  �&  �
i	  ��  �
  0U  �
�  @>  �
#  @  ��  `�  ��   f  ��  $�  ��  (P  ��  ,)x �	y   0)y �y   4�  �	y   8  �y   <F  �	y   @   �  -   �   �  -    
�  �  ��  *4�	�  'x �	y    'y �y   �  �	y     �y   �  �4   �  �4   �  �	y   �  �	y   �  �	y    L  �	y   $�  �	y   (H  �	y   ,�  ��  0 
�  #  �   2��F  �  �
�   )x �	y    )y �y   �  �	y     �y     ��  T  �	y   ��  �
�  �|  �	y   �  �	y   � �  ��  2ѣ  'x �	y    'y �y   �  �y     �y   'url �
�  |  �	y    �  �R  2���  'url �
�   �   �
�   ?  �	y   �   �4   �	  �	y   � �  ��  �    -    3  �  @% 3�  �y   (% 2��  'url �
�   �   �
�   ~  �	y   �?  �	y   ��  �	y   � �  �7  �  �  -    3�  ��  � 3�  �y   � 3�  �y   d�  +�  ��  @�   �  ,-   � +  ��  ��  +?  �y   ��  +�  ��   �  +  �i	  ��  +�  �y   ��  �  X  ,-    f  G  �5 	  y   �5   �  �5 F  �  ,-   � H	  �  �} r  y   �} �  �  -   � �  
�  �I F  y   `I �    -   _ y  �  ��   y   �� ND	a  Ourl 
�   <�   
i	   <   4   @ =V  +  a  |  -    �  l  �� ]  y   `�    y   x� P  y   t� m  y   p� �   y   l� 2  #y   `  $y   c	  *�   �    ]�  `�  P-   �j     �  s  �  �  D  �  k  A    =U  �$  z  �j  h� �  ��  d� �  �y   `�   �  ,-   � �  ��  `� �  �y   D� O   �y   @� >�  �#	  Lz  �  ��  #api �'(	  � "win �L         4  ��  @� -�z  b   a  "i �y   5   #    -�z  '   y  i �y    $�0  7{     �1  �   �     1  �   �      �  �  -    5�  ��r  W  ��  #mx �y   � #my �y   �#btn �#y   �?  �y   ?)  �y   (�  w  �  �y   �   �   �  �y   �   �   -dt  H   d  "i �y   �   �     �t  �    yw  �    (�  `  |  �y   �   �   �  �y   F  (  �  �y       �  "i �y   C  7    "lr ��  �  {  �  �y       �  �y   v  f      ��  ��{!  ��  ��} 3  u    1  ��  +3  ?  7  O3  �  x  C3  �  �  73  .  $  1  [3  ��}g3  N  �  l3  h  d  x3  �  �  �3  �  �  �3  �  �   �3  Zu   ]  �=  �3  �  �  4  0  &  4  {  m  ]  4  �  �  +4  �  �  74  �  �    �3  �  U  �3  �3   &�3  �u  �   �3  0  *  �3  T  N  �3  r  p  &�3  .v     �3  ~  |      �2  �v   �  �J  �2  �  �  �2  �  �  �2  �  �  �2  �  �2      �2  �  �2  V  @  �2  �  �2  ��{�2  �  �   3  �  3  �  �        8w  !"   wx  k        �s  !"   �t  !!   �w  !   ex  �    
�  5  �
4!  H  ��  #x �
y   � #y �
y   �#w �
!y   �#h �
(y   �  �
	y   ;	  7	  �  �
	y   P	  L	  �  �
	y   k	  c	  )  �
	y   �	  �	  |  &	y   �	  �	  P  '	y   �	  �	  �  (	y   
  
    -	y   E
  ?
  �  .	y   f
  ^
  (i   �  "i �
y   �
  �
  ~   �  �
4   �   �
�  ��}�  �
y   �
  �
  �  �
y   �
  �
    -�$  /     M  y   �
  �
   (�   ^  "i 1y     	  �   "box 2�  M  G    3y   �  �  x  4y   0  +   �   <�  o  �  �  c  �  �  Y  �  �  O  �  �  E  �  �  .;  @O+  u�} �  �&    �&  �   ER    �  �           +  )  �  8  4  �  M  I  �  c  _  �  v  t  .�  $  �  ~   @�&  u�}  (�   F  "i Ly   �  �  �   "run M�  �  �    Ny   *  "  x  Oy   �  Sy   Y  G  o  Wy     �  �  `4   Q  G    b�  ��}	  cy   �  y  R  gy   �  �  Q�)  8     sy   �  �     �   ;  y   �  �  -�'     w  i �y    �   �  �y   #    �  �y   �  ~       �  -    
�  
F  �  �
0  x �
y   y �
$y   w �
+y   h �
2y   �  �
9y   �  �
Ky   �  �
"4   �  �
4y   bw �
	y    3  �
|  x �
#y   y �
*y   w �
1y   h �
8y   �  �
?y   �  �
P4    5.  g
p  �  ��  #key g
y   � len h
	y   -�p  Y   �  "i �
y     �      pp   pp  P   p
  %   %  #  &1   �p     2   7  /    A>   pq   �  �
AE   �q   �  |
Rd   �q   �q  $   t
L   �q   �q  <   x
p  W   y  u   �  Dr   Dr  b   �
�  �  �  �     �  �  &   dr  "      �  �    S�p  �b  �  8K!  @�   �p  �    Mq  �    �  U
   c U
%  len V
	y   i Y
y     �  >
>   len ?
	y   i B
y     9�   9
9�  4
b   ,
d   len -
	y    9)	  %
5i  
�r  8   ��   #url 
#V  �  �r  �    �r  !"   T  
�   �  
y     
�     
�  Ur  �	�m  �   �:�   �	�m  5   �!   �m  !"   :b  �	hm  V   �!!   �m  !"   :|  �	m  O   �@!   `m  !"   �  �	r!  O  �	"V  url �	
�  �  �	�    �  �	�!  �  �	�  src �	-V   !*  �	y   �!  O  �	V   3  �	"  src �	$V  dst �	/�  !	  �	8y   i �		y   j �	y   c �	  hex �	"       !"  -    >�  N	y   DX  �  �u'  #url N	V  �   U	�       �  q		y   P  J  �6  �X   �X  S   U	�"  �6  r  p  &�6  �X  S   �6    }    �0  6Y   6Y  .   j	�"  1  �  �  1  �  �   u'  �Y   �  x		�&  �'  �  �  �'  	  �  �  �'  �  R  �'  �  k  �'    �  �'  �  �  �'    �  �'  �  �  �'    �  �'  �  �  �'  �  \   (  (  \  J  (  ��}$(  ��~0(  �  �  <(  �  �$  A(  �  x  M(  �  �  Y(  +    e(  {  m  q(  �  �  }(  *  z$  ~(    �  �(  U  �(  �  �  �(  �  �  �(  �  �  &�(  d  �   �(    
     $`*  �Z   y  #|*  A  ?  p*  M  K  y  �*  [  Y     �(  �  p&  �(  u  e  /Z)  i^    %  _)  �  �  k)  �  �  w)    	   �(  �  �%  �(  '    �(  �  x  �(  �  �  �(  	    )      )  &  $  )  �  �%   )  3  1   -)  �  .)  C  ?  :)  X  V    /�)  �e  �   �%  �)  f  b   /�)   g  �   &  �)  �  �  	�g  �)  Ps R��}��}"2Q��}2  /�)  �g  �   X&  �)  �  �  	ah  �)  Ps R��}��}"4Q��}2  H)  
  M)          &�)  �f  *   �)  �)  S   M   	�f  �)  Ps Qw     W6  �_      ~		7'  s6     y   6  �   �   �6  �   �   g6  !  �     �6  ,!  "!  �6  f!  \!  �6  �!  �!  �6  /  �6  �!  �!     ?6  �d   �d  M   W		_'  J6  �!  �!   	�Y  xa  8�*  ��    m  ��)  �  �y   �  �/y   y 	y   x 	y     	y   m  	y   �  	y     		y   �  
	y   2  	y   �  	y   �  	�)  �  	y   �   	�)    	�)  �  �  �(  �  �  len y   +  y   �  y     #y   i )y   run ,%�  �  -y   �  D%�  lr K0�      �)  E  fy   H)    yy   �  zy   �  �y   &  �y     �y   �  �y   -)  �  ~y    �  �y   n   �y     Z)  run �!�   �)  run �!�  *  �y   �  �y    �)  run �!�   �)  run �!�   run �!�    ^  	!y   �  	!y     y   �)  -    V.  �d  _  �`*  0�  �%�  "  �!  6x �/y   �"  �"  6y �6y   r#  `#  B�  =y   � B  Hy   �"box ��  %$  $   !�  �y   �*  �  �#V    �-y   len �	y    >  (+  D  ($V  �   -
i	  �  .	y   �  /
+  '   0	y   \  1
+  R  2	y   p 4V  c 6      +  ,-   �   -+  ,-   � �  ��+  �  �%V  len �/y   ;  	y   �  �  x+  i y    �  "y     �  ��+  �   �(V  <  ��  �  ��   WR	  ��N  D  �R/  0�   �*V  n$  `$  0�  �:�  �$  �$  0'   �Ey   @%  2%  <  ��  �%  �%  �  ��  �%  �%  �  ��  Q&  3&  (�  �.  [  ��  �  �y   �&  �&  �  ��  ��}(<  �,  m  �  N'  H'  �  ��  p'  l'  �  �y   �'  �'   (-  �,  �  ��  �  �y   �'  �'   �1  �T   K  �Q-  �1  �'  �'  �1  (  (  K  �1  �1  �1  	U  �E  Pv Rw s "#�   �P  �5  m-  Ps R��{ �P  �5  �-  Ps R��{ �P  �5  �-  Ps R
��{����" Q  �5  �-  Ps R
��{]���" "Q  �5  �-  Ps R
��{����" BQ  �5  .  Ps R
��{����" bQ  �5  3.  Ps R
��{����" �Q  �5  U.  Ps R
��{����" �R  �5  r.  Ps RN�   	�T  �5  Pv R_�    �0  &O   &O  p   ��.  1  (  (  1  (  (   �0  �Q   Z  �/  �0  7(  3(  �0  R(  N(  $�0  �Q    i  |�0  q(  m(  �0  �(  �(    O  |1  3/  Ps  	�O  %1  Pv R��{Qs   Z  ��0  D  �0V  I  �	y   p �V  g0  �  �y   �   �#  3  �y   �  �+  '   �y   X0  <   �  �  
!�  �  %V  [  )V  �  !y   �  "�  :0  m   *  �  !1V  �  #)y    �  )1V  �  +)y        <  W �    �  eV  R  gy   6  m�     �  ��0  R   �0V  p �V  m  �  �  �+  �  �y     �   |�0  �  |*�    |>�   !�  t�  %1  A  t4!  �  v�   C	  ]�  d   �  �|1  0<  ]5�  5)  �(  0�  ]L�  i,  a,    ^�  �,  �,   !1  #�  �1  tag #4V     (�2  �  (,V    (D�2  p +V  �  ,
i	  �  ,�  �  2y   �  <y   ,2    n�2  v  o�2  cnt py   vp qV   U2    ��2  cnt �y   vp �V   f2  vp �V   w2  vp �V   vp V     
�  y   �2  -    !�  �y   3  url �0V  �  �;�  !	  �Jy   �  �V  i y   hex 	3  val 
y   j "y           3  -    c  ��3  _  �%V  �  �;V  �  �O�  !	  �]y   >  �
�  �3    �V  �  �y   �  �y   �   �y    �3  �  �y   �   �y      �V  �  �y   �   �y   �  �y      6  �D4  url �(V  >  �3�  !	  �?y     �V  �  �V  k  �	y    !�  xy   a4  �  x'V   !\  py   ~4  �  p'V   !�   iy   �4  �  i(V   !r  ]y   �4  �  ])V   !  Ry   �4  �  R*V   !?  Hy   �4  �  H.V   !&  @y   5  �  @-V   !�  3y   ,5  �  3+V   !G  y   U5  Y   #V  �  !	y    !�  �y   �5  �  �$V  �5  len �y   �  �4   i �y   c �     p �V  r �y   g �y   b �y     CV  �y       c   �?6  6s1 �$V  �,  �,  6s2 �4V  �,  �,     "c1 �  -  -  "c2 �  !-  -    �  �W6  �  �)�    !n  ��   �6  url �,V  �   �=V  "  �-V  len �:y   -  �	y   �  �4   �  ��   i �y     !,  ��   �6  url �-V  i �y     4U5  �  +  �<  e5  B-  ,-  �5     S7  �5  �-  �-  �5  �-  �-  �5  �-  �-  �5  .  �-   q5  (   �7  v5  ".  .  �5  >.  8.  �5  3   �5  a.  U.  �5  C   �5  �.  �.     �  �5  �7  Ps R��   �  �5  �7  Ps R �   �  �5   8  Ps R�   �  �5  8  Ps R�   �  �5  :8  Ps R��     �5  W8  Ps R��     �5  t8  Ps R��   +  �5  �8  Ps R�   @  �5  �8  Ps R�   U  �5  �8  Ps R��   j  �5  �8  Ps R��     �5  9  Ps R�   �  �5  "9  Ps R$�   �  �5  ?9  Ps R+�   �  �5  \9  Ps R1�   �  �5  y9  Ps R6�   �  �5  �9  Ps R;�   �  �5  �9  Ps R@�     �5  �9  Ps RE�   '  �5  �9  Ps RM�   <  �5  
:  Ps RT�   Q  �5  ':  Ps R[�   f  �5  D:  Ps R`�   {  �5  a:  Ps Rf�   �  �5  ~:  Ps Rl�   �  �5  �:  Ps Rt�   �  �5  �:  Ps Ry�   �  �5  �:  Ps R��   �  �5  �:  Ps R��   �  �5  ;  Ps R��     �5  ,;  Ps R��   #  �5  I;  Ps R��   8  �5  f;  Ps R��   M  �5  �;  Ps R��   b  �5  �;  Ps R��   w  �5  �;  Ps R��   �  �5  �;  Ps R��   �  �5  �;  Ps R��   	�  �5  Ps R��    1,5  �  p   �?<  <5  /  �.  H5  /  /   1,5  `     �|<  <5  @/  8/  H5  Xk  <  P	�� &�-�   15  p    ��=  5  {/  o/  5  �    S   3j=  5  �/  �/  �  �5  �<  Ps R��   �  �5  �<  Ps R�   �  �5  =  Ps R�   �  �5  3=  Ps R�     �5  P=  Ps R�   	  �5  Ps R �    �  �5  �=  Ps R��   �  �5  �=  Ps R��   	�  �5  Ps R��    1|1  x  �  �SD  �1  �/  �/  |1  �    ^   #�C  �1  30  /0  �  �5  >  Ps R,�   �  �5  ;>  Ps R2�     �5  X>  Ps R6�     �5  u>  Ps R$�   +  �5  �>  Ps R;�   @  �5  �>  Ps R>�   U  �5  �>  Ps RA�   j  �5  �>  Ps RD�     �5  ?  Ps RG�   �  �5  #?  Ps RJ�   �  �5  @?  Ps RM�   �  �5  ]?  Ps RP�   �  �5  z?  Ps R��   �  �5  �?  Ps RS�   �  �5  �?  Ps RW�     �5  �?  Ps RZ�   '  �5  �?  Ps R]�   <  �5  @  Ps R`�   Q  �5  (@  Ps Rf�   f  �5  E@  Ps Ri�   {  �5  b@  Ps R-�   �  �5  @  Ps Rl�   �  �5  �@  Ps Rr�   �  �5  �@  Ps Rx�   �  �5  �@  Ps R}�   �  �5  �@  Ps R��   �  �5  A  Ps R��     �5  -A  Ps R��   #  �5  JA  Ps R@�   8  �5  gA  Ps R��   M  �5  �A  Ps R��   b  �5  �A  Ps R��   w  �5  �A  Ps R��   �  �5  �A  Ps R��   �  �5  �A  Ps R��   �  �5  B  Ps R��   �  �5  2B  Ps Rb�   �  �5  OB  Ps R��   �  �5  lB  Ps R��   
  �5  �B  Ps R��     �5  �B  Ps R��   4  �5  �B  Ps R��   I  �5  �B  Ps R��   ^  �5  �B  Ps R��   s  �5  C  Ps R��   �  �5  7C  Ps R��   �  �5  TC  Ps R��   �  �5  qC  Ps R��   �  �5  �C  Ps R��   �  �5  �C  Ps R�   �  �5  �C  Ps R�     �5  �C  Ps R�   	  �5  Ps R�    �  �5  D  Ps R'�   �  �5  9D  Ps Rm�   	�  �5  Ps Rs�    4-+  |,  �  ��E  8+  J0  B0  D+  w0  i0  P+  \+  $-+  �,    �   �D+  �0  �0  8+  �0  �0  �   P+  1  1  \+  ,1  &1  /h+  �,     �D  m+  F1  D1   �0  �,   �,  `   )E  1  Q1  O1  1  ^1  Z1   �0  �-   �   �E  �0  r1  n1  �0  �1  �1  $�0  �-   �   |�0  �1  �1  �0  �1  �1    &x+  �-  '   y+  �1  �1      4�1  T.  �  ��[  �1  �1  �1  �1  �1  �1  �1  
2  2  �1  ��~�1  ��~�1  
  �1  %2  !2  �1  <2  42  U5  /     FIF  e5  a2  [2  	0/  �6  P��~  U5  }/   &  K~F  e5  �2  }2  	�/  �6  P��~  ,5  �/   �/     M �F  <5  �2  �2  H5  	0  <  P��~  ,5  �1   �1     b&�F  <5  �2  �2  H5  	�1  <  Pw   ,5  K2   K2     e)6G  <5  �2  �2  H5  	\2  <  Pw   ,5  �2   �2     h'sG  <5  �2  �2  H5  	�2  <  Pw   ,5  Z3   Z3     �"�G  <5  �2  �2  H5  	p3  <  P��~  ,5  �3   �3     �%�G  <5  3  3  H5  	�3  <  P��~  ,5  �3   �3     �#-H  <5  )3  #3  H5  	�3  <  P��~  ,5  �3   �3     �$kH  <5  K3  E3  H5  		4  <  P��~  ,5  =4   =4     �$�H  <5  m3  g3  H5  	S4  <  P��~  ,5  p4   p4     �#�H  <5  �3  �3  H5  	�4  <  P��~  ,2  1  (I  12  ��~=2  �3  �3  I2  4  �3  	5  ,5  Pw   U5  ;5   F  �#]I  e5  24  *4  	Q5  �6  P��~  U2  Q  �I  Z2  b4  X4  U5  �9   �9     �'�I  e5  �4  �4  	�9  �6  Pw   38  ,5  �I  Pw  	
9  5  Pw   ,5  �5   �5     �!J  <5  �4  �4  H5  	�5  <  P��~  �1  p  xJ  �1  ��~2  ��~2  �4  �4   2  �4  �4  S6  �5  gJ  Pw R��} 	P7  ,5  Pw   ,5  �6   �6     k(�J  <5  5  5  H5  	�6  <  Pw   ,5  �7   �7     �#�J  <5  5  5  H5  	8  <  P��~  ,5  8   8     �$1K  <5  ?5  95  H5  	�8  <  P��~  ,5  �8   �8     �"oK  <5  a5  [5  H5  	�8  <  P��~  ,5  >9   >9     �"�K  <5  �5  }5  H5  	T9  <  P��~  a4  :   {  �AL  q4  �5  �5  2:  �5  �K  Pw R��   C:  �5  
L  Pw R��   T:  �5  'L  Pw R��   	e:  �5  Pw R��    D4  .;   �  ��L  T4  �5  �5  B;  �5  �L  Pw R�   S;  �5  �L  Pw R�   k;  �5  �L  Pw R �   �;  �5  �L  Pw R)�   	�;  �5  Pw R/�    ,5  �;   �;     �0M  <5  �5  �5  H5  	�;  <  P��~  �4  �;   �  �%�M  5  6  6  <  �5  pM  Pw R�   <  �5  �M  Pw RM�   4<  �5  �M  Pw RY�   	I<  �5  Pw R`�    �4  ~<   �  �&�N  �4  ,6  "6  �<  �5  N  Pw R�   �<  �5  !N  Pw R��   �<  �5  >N  Pw R��   �<  �5  [N  Pw R��   �<  �5  xN  Pw R��   	�<  �5  Pw R��    �4  (=   �  �"}O  �4  _6  Y6  <=  �5  �N  Pw R��   S=  �5  �N  Pw R�   m=  �5  O  Pw R��   �=  �5  )O  Pw R��   �=  �5  FO  Pw R��   �=  �5  cO  Pw R��   	�=  �5  Pw R��    �4  �=   �  �!�P  �4  �6  z6  >  �5  �O  Pw R��   >  �5  �O  Pw R�   .>  �5  �O  Pw R��   C>  �5  P  Pw R��   X>  �5  1P  Pw R��   m>  �5  NP  Pw R��   �>  �5  kP  Pw R��   	�>  �5  Pw R��    ~4  �>   �>  G   �  Q  �4  �6  �6  �>  �5  �P  Pw R��   �>  �5  �P  Pw R��   	?  �5  Pw R��    ,5  (?   (?     � >Q  <5  �6  �6  H5  	>?  <  P��~  ,5  [?   [?     �"|Q  <5  �6  �6  H5  	q?  <  P��~  ,5  �?   �?     �&�Q  <5  �6  �6  H5  	�?  <  Pw   f2  �  (R  k2  7  �6  �A  ,5  �Q  Pw  B  ,5  �Q  Pw  ?B  �5  R  Pw R��} 	NB  ,5  Pw   ,5  �@   �@     fR  <5  27  ,7  H5  	�@  <  P��~  ,5  �@   �@     �R  <5  Z7  T7  H5  	�@  <  P��~  ,5  A   A     
�R  <5  �7  |7  H5  	A  <  P��~  ,5  9A   9A       S  <5  �7  �7  H5  	OA  <  P��~  ,5  lA   lA      ^S  <5  �7  �7  H5  	�A  <  P��~  w2  �  �S  x2  8  �7  U5  C   C     +�S  e5  D8  B8  		C  �6  Pw   �A  ,5  �S  Pw  !B  ,5  �S  Pw  	�B  ,5  Pw   /  �5  T  Pw RN�   y/  �5  #T  Pw RC�   �/  �5  @T  Pw RN�   �/  �5  ]T  Pw RC�   �/  �5  zT  Pw RT�   �/  �5  �T  Pw R_�   L0  �5  �T  Pw Ri�   d0  �5  �T  Pw Ru�   �0  �5  �T  Pw R~�   �0  �5  U  P��~R��   �0  �5  )U  Pw R��   1  �5  FU  Pw Rz�   <1  �5  cU  Pw R��   T1  �5  �U  Pw R��   u1  �5  �U  Pw R��   �1  �5  �U  Pw R��   �1  �5  �U  Pw R��   �1  �5  �U  Pw R��   2  �5  V  Pw R��   72  �5  .V  Pw R��   w2  �5  KV  Pw R��   �2  �5  hV  Pw R��   �2  �5  �V  Pw R��   �2  �5  �V  Pw R��   3  �5  �V  Pw R��   =3  �5  �V  Pw R��   V3  �5  �V  Pw R�   �3  �5  W  Pw R�   �3  �5  3W  Pw R�   �3  �5  PW  Pw R*�   "4  �5  mW  Pw R8�   94  �5  �W  Pw R@�   l4  �5  �W  Pw RN�   �4  �5  �W  Pw R[�   �4  5  �W  P��~ 75  �5  �W  Pw Rh�   t5  �5  X  Pw Ru�   �5  �5  0X  Pw R|�   �7  �5  MX  Pw R��   {8  �5  jX  Pw R��   �8  �5  �X  Pw R��   :9  �5  �X  Pw R��   �9  �5  �X  Pw R��   �9  �5  �X  Pw R��   �9  �5  �X  Pw R2�   :  �5  Y  Pw R��   �:  �5  5Y  Pw R��   �:  �5  RY  Pw R��   �:  �5  oY  Pw R��   ;  �5  �Y  Pw R��   &;  �5  �Y  Pw R�   �;  �5  �Y  Pw R6�   �;  �5  �Y  Pw R>�   r<  �5   Z  Pw Ro�    =  �5  Z  Pw R��   �=  �5  :Z  Pw R��   �>  �5  WZ  Pw R��   $?  �5  tZ  Pw R�   W?  �5  �Z  Pw R�   �?  �5  �Z  Pw R�   �?  �5  �Z  Pw R��   �?  �5  �Z  Pw R��   @  �5  [  Pw R��   i@  �5  ![  Pw R��} �@  �5  >[  Pw R"�   �@  �5  [[  Pw R*�   A  �5  x[  Pw R��   5A  �5  �[  Pw R&�   hA  �5  �[  Pw R0�   	�A  �5  Pw R:�     4�0  C    ��`  �0  l8  N8  7�0  `� ��0  )  �0  9  9  �0  ��_�0  W9  G9  $R/  D   8  �]/  �9  �9  8  i/  :  :  u/  `:  ":  /  \  `  �/  �;  �;  �/  ��Y�/  �;  �;  �/  ��[�/  <  	<  �/  �  �_  �/  O<  E<  �/  �  �_  �/  �<  �<  �0  H   �  
(]  1  �<  �<  �  1  �<  �<    �/  �  �/  �<  �<  �/    T_  �/  �/  �=  ~=  0  ��Y:0  4  r]  ;0  G0  �=  �=   /0  �L  M   �]  0  >  >  !0  />  ->  -0  ?>  9>   �1  �M   C  F!^  �1  d>  b>  �1  x>  v>  C  �1  �1  �1  	�M  �E  Pu Rs w "#�   �I  �5  /^  Ps R
��W����" �I  �5  Q^  Ps R
��W����" �I  �5  s^  Ps R
��W����" �I  �5  �^  Ps R
��W]���" �I  �5  �^  Ps R
��W����" J  �5  �^  Ps R
��W����" 8J  �5  �^  Ps R
��W����" XJ  �5  _  Ps R
��W����" 	L  �5  :_  Ps RN�   	�M  �5  Pu R_�    �0  �J    R  M�_  �0  �>  �>  �0  �>  �>  $�0  �J    a  |�0  �>  �>  �0  �>  �>    	�H  %1  Pv Rw    	 H  |1  Pv   X0  p  Y0  �>  �>  	�G  |1  P��Y   g0    h0  t0  	?  �>  �0  �  �0  Q?  M?  �0  E   E  m   m)j`  1  f?  d?  1  s?  q?   $�0  F   �  y�0  ?  }?  �0  �?  �?  $�0  F   �  |�0  �?  �?  �0  �?  �?          1�+   N  �   �xa  �+  �?  �?  �+  z@  t@  �+  �+  DN    �  �Na  �+  �@  �@  �  �+  �+  �@  �@  	ZN  �5  PsRv    5N  |1  ba  Pv  	�N  �[  8�0  `�   1�*   U  "  ��b  �*  ��[�*  �@  �@  �*  ��[�*  \A  LA  �*  ��_�*  �A  �A  �*  "B  B  7�*  ��  ��*  x  �b  �*  �B  �B  �U  -+  b  P��_Ru  �W  �+  @b  P��[R��[Q��[ �W  �+  Vb  P��[ �W  �+  zb  P��[R��[Q��[ 	�W  �+  P��[  	6W  -+  P��_Ru   4@!  j  �  ��c  W!  ��{7K!  @� ��!  Hj   E  �		�b  �!  �C  �C   c!  T  �c  d!  ��}Y�!  c  �		qc  .�!  .�!  .�!  c  �!  D  �C  �!  xD  hD  �!  y  �!  �D  �D  "  �  "  ��{    $r!  �l   �  �		�!  �D  �D  }!  E  E    r!  l   l     �	�c  �!  )E  %E  }!  EE  AE    �j  !"   Z�   �n  s  �7�   � $�   �n    �  
�   ^E  XE  &�   �o  �   �   �E  |E  [�6  �o  1   
$\d  .�6  &�6  �o  1   �6    ?6  �o   �o  O   
�d  J6  �E  �E    �o  !"      �   d  4|	  r       0}    [  �  2   �  R  E   5q	  	S   X   r   r   r   r   r    6int !  
�   �   �   r    �  �   �   �   r   r   r    h  �   �   �   r   r    0   �      I  #   
    2    �  7  
  ,  2     ]  �  
]   �  4m  �  	r   � 
  m  2    
�   }  2    �  ,  �	D  �  T   F  o    �  �  �    �  1   �  �  !�  E  "�  �  %   �  &  $�  '!  (�  (:  ,r  )�  07   *�  4�  +�  87  .g  <-  /�  @�  0�  D�  1�  Hn  2�  L�  3  P[  45  Tz  5Y  X@  8s  \�  9�  `�  :�  d�  ;�  h*  <�  l�   =�  p�  >�  t   ?  x*  @�  |7  A,  �Y  B@  ��  CU  ��  F_  ��   G_  �  H_  ��  I~  ��  J_  �  M  �E  N�  �h  O�  �  P�  �  Q�  ��  R
  ��  S7  �K  TZ  �1   Un  ��  V�  ��  W  �   X  ��  [�  � O  O     D  E   h  h   �  Y  E   �  E   h   t  �  E    �  8�  r   �  O   �  r   �  O  O   �  �  �  r      �  r     O  �  r    �  r   !  O  E   r      r   :  O  r    &  9   g  O  r   r   G   y   �    ?  �  r   r   r   r   r    l  �  r   r   O  r    �  �  r   r   O  r   r    �  �  r   r   O   �    r   r   r   r   O   �  5  r   r   r   r   r   r      T  9   T  r   �    }  :  s  E   r   h   ^  �  E   �  h   �  9x  �  �  O   �  �  �  O  h   �  r   �  O  O  h   �  �  �  O  r    �  �    O  O   �  r   ,  �  O  :   h  @  O   1  U  r   �   E  ;&   Z  y  y  y  y   r   d  r   �  r   r   r    �  r   �  r   �  r    �  r   �  r   �  h  r   �  r    �  r   
  r   �  h  r    �  r   7  r   E   h  r   E   y     r   Z  r   E   h  r    <  r   n  r    _  r   �  �  �  �   s    ]�  �  �  T  0-�  �  .�      /r   (M  0r   , 
  �  2   '  �	  ~  	r    W  	r   �   
  K  
�	  (F   
�	  ��  !
�	  ��  $	r   �/  %	r   �  (�  �]  1�	  �<f  2	r   � 
  �	  2    
  �	  2   ? 
  �	  2    
�  �	  2   ? �  3�  =�  6�	  �  �  �  �  �  �  �  &   >sys �  `N $2	I
  &id 3    4�    :  5)
  
I
  e
  2    �  7U
   H C  8r   �G 
}  �
  2    /  :�
  `J 	  ;r   DJ  >�
  &key ?  �  @
�
    
  �
  2   �   A�
  
�
    2    �  C�
  �> >  Dr   �> ?�	  O�1    �r   ��  �   ��  key �r   � �  }  len �r   �E  �E   ߔ  �    r  fr   ��  �  ��  	�  fr   � 	�  f$r   �mx f/r   �my f7r   �x i	r   �E  �E  y j	r   \F  TF  �  u	r   �F  �F  �  v	r   �F  �F  fy �	r   �F  �F  �  }  idx zr   �F  �F  �  {r   G  G  Z�  �  ��  �   !�  ֒  �  i�  �  DG  @G   !�  �  �  j�  �  \G  ZG   6�  #   @�  Er   ��  %   �  mx E r   � my E(r   �btn E0r   �  P  �r   �  �  ��  	e  �r   � 	�  �%r   �	�  �0r   �	�  �;r   �x �	r   wG  kG  y �	r   �G  �G  �  	r   H  H  �  	r   >H  :H    	r   UH  QH  A�  	r   fy 0	r   nH  fH  "�  �   S  i r   �H  �H  �  idx r   �H  �H  iy  r   �H  �H  8  (O  I  I  \�  ^    !�  %�  �  �v  �   I  I   '�  =�  �  ��  1I  /I    (�  �D�  �  ��  �  �
�	  ��~len �	r   HI  @I  ��  �   #�  �ȋ  {   �#  	�  �'O  � len �	r   gI  eI  B7�  w <�     C�  �=  )len �r    DW  �Ċ  \   ��  �   �!O  sI  oI  �  �4O  �I  �I  	�  �KO  �	�  �eO  �cb �~�  ��  �   #  ��  �   �  	�   �!O  � 	�  �4O  �	�  �KO  �cb �d�  ���     Ea  ���  V   �(�  [��  3  ��  F@d�  �  e�   M  f&   (0  g&   ,[  h�	  0*uid i�	  1�  j�	  2*gid k�	  3�  l�  4 G#  m4  �  o	r   �I  �I  �  p�  �I  �I  �  �  u	r   �I  �I  b  i wr   #J  J  m     {r   QJ  KJ  �  �r   oJ  kJ  x  i  �  �r   �J  �J  �  �r   �J  �J   ��  F   idx �r   �J  �J      
&   �  2    +�  HD�  :   �^    H&
  �J  �J  �  H8O  �J  �J  x HBr   �J  �J  y HIr   K  K  dw HPr   �dh HXr   �cx H`r   �cy Hhr   �cw Hpr   � ch Hxr   �$,{�  -��  +k  E�  :   ��  �  E
  #K  K  �  E2O  >K  4K  x E<r   kK  eK  y ECr   �K  �K  	�  EJr   �	�  EUr   �,?�  -��  #p  "Ć  D   �  	�  "E   �  $�  �r   0�  �  �o  U  �$O  Vf  
�	  ��~)len r   �  
�  VM  	r   P $�  �O  ��  v   ��  key �'O  � ʄ  O   i �r   �K  �K    %  �`�  �  �2  xml �$�  � ptr ��  �K  �K  ,  �  ��  �K  �K  z  ��  L   L  <    |  �r   "L  L  i �r   FL  @L  �  ��  bL  ^L    ��  vL  rL  L    �  ��  �L  �L  �  �r   �L  �L  =  ��  �L  �L  �  ��  M  M  "��  H   �  k �r   LM  HM   "@�  L   �  k �r   `M  \M   ہ  �  �  �  3�  �   ��  �   �  �  
�  �    %q  ���  �  �j  buf ��  rM  pM  ptr ��  M  {M  W  �  ��  �M  �M  &  ��  �M  �M  B  ��  �M  �M    �  �@  �r   �M  �M  r  ��  �M  �M  �  ��  �M  �M    ��  N  N  �  �r   N  N  Z�  �  q�  �  ��  �  ��  j  Ƀ  �  ��  �  ��  �  h�  j  ��  �    He  �(�  8   ��  I�  ��  pN  fN  src �+O  �N  �N  n �4r   �N  �N  i �	r   �N  �N   J/  m�  .�  m!r   .y  m/r   Kid }O   /H  c   |   �2  id c'O  � !  i dr   O  O    %W  \�~  N   �c  I  \!O  �   \3�  � /  H ~  �   ��  api H�  0O  *O  �  Ir   @J  0�  &�   ~     ��  s &O  MO  IO  c &$r   aO  ]O   $�  �  h}  �   �X  �  O  � (  3O  �R  	r   uO  qO  �  	r   �O  �O  �}  8   i  r   �O  �O  �}  X    0�  r   0}  5   ��  s1 �  � s2 +�  �n =h  �p1 O  �O  �O  p2 O  �O  �O  6}  &   i h  �O  �O    L�  r   �  Mval !r    N�  �  �   �z  1�  � 1�  �2�  �O  �O  O�  �   �     mg  �  ?P  ;P  �  QP  OP  3�  �  �   �  �  �  �   P#   �  �   �31  '#  S�   �  ��  21  iP  [P  ��        %Q   �
  N|	  �       D�  [B  �k   �   �    @    �   �   �   �  Oint  �   �   �  B-   �   T   �  �  �  S  �  �  &  C   @   x   q  %�   Co  3  A  4�    ;  5  �  6	\    �  &  C  HAI  �  Bh   b  C	\   @�  D�  D u  'U  PJ  �J}  K  Kx     L	\   � Q )	�  '�  *	\   '�  +	\   '  ,
�  '  -�  'M  .�  'i  /	\   '�  0   �  �  -   �  �  R�    I  S    =\   =   �     �  K  1}  DD<L  Ekey =
L   �  >  @ �  \  -   ? [  ?*  \  x  -      �  -    DHR�  �  S
L   �  T  @1  U	\   D �  V�  2P[  �  \
L   �  ]  @  ^
#  D  _	\   DG  `	\   H�  a  L �  �  9  -   -      b�  2	g�  �  h�   �  i�  �  j	\   	�  k	\   	K  l  	 9  �  �  -    �  mE  T$� r	�  �  t�   �  u	\      �  x�    �  y	\   $ `  |�  $ �  }	\   N �  ��  N �  �	\   �    ��  � {  �	\   � |  �
�  � �  �	\   �   ��  � �  ��  �   �   �  4   �  F-   �� �  �  -    9  �  -    �  �  -    �   �  -   � UV�  =�   �  �  �  ��  �  $  -    �  4  -    B-   %p  �   3  �  �  7  �  �     f  .4  20�  A  1p   �  2
�  �  3	\   �  4	\   �  5	\    �  6|  �  �  -    .�  9�   �  �    -   " .1  A�  ��  28L�    M�   Epos N	\     O	\   �  P	\   �  Q	\   �  R�    S�  $  T	\   4   U  2@Z�  �  [�   �  \�  81  ]	\   <�  ^
�  @   V  _�  /�  �<�  c   ��  �  �'�  � 	8  �  �P  �P  	  �  �P  �P  	>  �  �P  �P  V�  �F  g�  R	  o�  �F  ��  R	  ��  �F  ��  R	   6'  �  �  n  �'\   P  �:   7&  �  �  n  �&\   P  �9   6�  �  �  n  �!\   P  �4   �  �  �     �;  n  �.\   � P  �A  ��  �E   6�  �  c  n  �+\   P  �>   7i  �  �  n  �,\   P  �?   6s  �  �  n  �!\   P  �4   7�  �  �  n  �"\   P  �5   7�  �  	  n  � \   P  �3   /�  xT�     �(	  �  x"�  �  x  t�  H�  
   �R	  �  t'�  �  /�  dT�  �   �
  (�  d!�  �P  �P  �  d5�  ��  dG  �
  �	  i e\   Q  Q  D  ��      f3D  >Q  6Q  )D  aQ  [Q    �I  ʭ    (  m	�I  {Q  wQ  �I  �Q  �Q    =  ^  �  k   ��
  �  ^(�  � �  ^<�  �var _�
  �Q  �Q  <<  �   �  _X<  �Q  �Q  L<  �Q  �Q  "d<  �  e<  �Q  �Q  D  �   �  �3D  R  R  )D  0R  (R      �  C  P\   \�  �   �i  (�  P%�  QR  MR  (�  P9�  gR  aR  #fn Q&  �	  T�  �R  R  �I  ��    ��     U�I  �R  �R  �I  �R  �R      >  ��    ��  �  >"�  � 9  >6�  �>�  ?�  ��y	�  F  �R  �R  HE  -�   -�  J   D*  ]E  �R  �R  RE  �R  �R  3�I  ?�   ?�     ��I  �R  �R  J  CS  ?S    �<  ��   �  Hf  �<  [S  WS  ��  �<  Pv R��w  ��  I  ��  =  P��w  /�  :@�     �  �  :�  � �I  @�   @�     ;W�I  $� X�I   �I  tS  rS  �I  S  }S  8�I  @�     �I  �S  �S     	  1\    �     �;  �  1"�  � #arr 16  � >  #  ̫  Q   ��  �  #'�  � #arr #;  ��  #D\   �	M  (�  �S  �S  �  I   /�  ��  0   ��  �  !�  � #arr 5  ��  F  �	M  �  �S  �S   �    �  �   ��  �  (�  � #obj <  �#key M�  �  
�  
�  �  i \   T  �S  D  .�    �  3D  +T  #T  )D  NT  HT    j�  I   /�  ��  �   �q  �  �!�  � #obj �5  �#key �F�  ��  �W  �  ��  
�  C  i �\   nT  dT  D  :�    �  �3D  �T  �T  )D  �T  �T    �I  |�    �  �	�I  �T  �T  �I  �T  �T    �  �  P�  �   ��  �  �(�  � �  �<  ���  qH  ��  qH  ȩ  qH  ٩  �E   �  �  T�  �   �o  �  �'�  � �  �;  �
�  S  num �\   �T  �T  p ��  U  U  neg �\   3U  -U  '�  H   ��  H  ��  H  Ũ  �E   �  �  �  l  �=  �  �'�  � �  �;  �
}    9buf �$  �@n �\   XU  LU  i �\   �U  �U  )�  d     neg �\   �U  �U   ç  �G   '�  �G  G�  �G  g�  �G  ��  �G  ٧  �E   ?g  u  �  �  ��  (�  u.�  V  �U  	�  v�  4V  ,V  tok w�  eV  [V  	�  �  �V  �V  
S  l  	�  |  �V  �V  q<  ��   g  {	"  <  W  W  q<  w�   w�      �<  W  W  ��  �<  Pv Ru    �<  ��   t  }\  �<  )W  %W  ��  �<  Pv Ru   D  �  ~.�  3D  >W  :W  )D  TW  RW   �<  �   �  "   ��  �<  ^W  \W  -�  �<  Pv Ru   D  n�  0   �*�  3D  jW  fW  )D  �W  ~W   q<  ��   �  �R  <  �W  �W  q<  ��   ��     �<  �W  �W  ��  �<  Pv Ru    ��  I  �  =  Pu   �<  +�   =  w�  �<  �W  �W  ��  �<  Pv Ru   �<  I�   H  ��  �<  �W  �W  ��  �<  Pv Ru   D  w�    w�  '   z&  3D  �W  �W  )D  X  �W   D  �    �  2   �&J  3D  X  X  )D  4X  2X   q<  N�   �  �	�  <  AX  =X  q<  ��   ��     �<  VX  TX  ��  �<  Pv Ru    F�  �  Pu   �  �  �  ?�  A  ��  T  ��  (�  A/�  hX  `X  	�  B�  �X  �X  	5	  D  �X  �X  tok F�  Y  Y  
+  9  op H�  OY  GY  )��  0   �  n   L  q<  ��   ��  0   K<  vY  rY    )��     �  n   R  Gq<  ��     Q0<  q<  ��   ��     �<  �Y  �Y  ��  �<  Pv Ru     
l  �  	n   \  �Y  �Y  q<  �   w  [p  <  �Y  �Y  q<  ��   ��      �<  �Y  �Y  ��  �<  Pv Ru    �<  \�   �  ^�  �<  �Y  �Y  ��  �<  Pv Ru   A�    �  Pu  X�  �K  R��}Q��}Y0;  u   
'  �  	�  d  �Y  �Y  
2  T  	]  h  �Y  �Y  	�  i\   Z  Z  W�  q<  C  Pu  ^�  �  Pu   !�  q<  h  Pu  (�  �  |  Pu  1�  �<  �  Pu  H�  D  R��    D  �   �  .   J�  3D  Z  Z  )D  +Z  %Z   D  ;  P  3D  GZ  CZ  )D  ZZ  VZ   D  x�     P!3  3D  kZ  iZ  )D  uZ  sZ   D  K  P5^  3D  Z  }Z  )D  �Z  �Z   D  V  PI�  3D  �Z  �Z  )D  �Z  �Z   D  a  V�  3D  �Z  �Z  )D  �Z  �Z   D  �  V �  3D  �Z  �Z  )D  �Z  �Z   D  �  V3
  3D  �Z  �Z  )D  �Z  �Z   D  �  VF5  3D  �Z  �Z  )D  �Z  �Z   D  �  W`  3D  �Z  �Z  )D  [  �Z   D  �  W �  3D  [  	[  )D  [  [   D  �  W4�  3D  [  [  )D  )[  '[   D  �  X�  3D  3[  1[  )D  =[  ;[   D  �  X!  3D  G[  E[  )D  Q[  O[   D  �  Y7  3D  [[  Y[  )D  e[  c[   D  �  Y b  3D  o[  m[  )D  y[  w[   D  �  Y3�  3D  �[  �[  )D  �[  �[   D    YG�  3D  �[  �[  )D  �[  �[   D    Z�  3D  �[  �[  )D  �[  �[   D    Z!  3D  �[  �[  )D  �[  �[   GD   �     b3D  �[  �[  )D  �[  �[    �<  ��      Fs  �<  �[  �[  ��  �<  Pv Ru   ��    Pu   !�  �    �  �2�  �  �F�  �  ��  tok ��  P  �  n  �	\     9�  val !\   p "�        -    Z#    @�  �  �;  (�  ,�  8\  �[  	�  �  �]  �]  tok �  h_  _  
�    >�  &L  ��~	�  *  �`  �`  )E�  Q   �  var 2$�
  !a  a  �I  _�    _�     3�I  9a  5a  �I  La  Ja    �I  �  '  �I  Za  Ta  �I  ~a  ta   q<  ��   �  (q  <  �a  �a  q<  ��   ��     �<  �a  �a  ��  �<  Pv Ru    �<  �   �  +�  �<  �a  �a  ��  �<  Pv Ru   D  r�  ,   ,2�  3D  �a  �a  )D  �a  �a   �  I  ��  q<  �  Pu  ��  �  Pu   
  F  	  @  b  b  	�  F  ?b  5b  	�  G\   kb  ib  ��  q<  a  Pu  ��  �  u  Pu  ��  �<  �  Pu  ��  I  ��  =  �  Pu  ��  �<  �  Pu  �  D  �  R��   �  q<  �  Pu  H5�  =  �  P��|H F�  D    R�   U�  q<  (  Pu  -�  =  <  Pu  @�  =   
�  �   	�  c\   xb  tb  	�  e  �b  �b  	�  f\   �b  �b  	�  g\   �b  �b  
�  f   	  k!  �b  �b  �  q\   D    m6�  3D  c  c  )D  c  c   �<  ��     l-   �<  4c  0c  ��  �<  Pv Ru   ��  =  A   Pu  ��  �  U   Pu  -�  q<  Pu   Z�  q<  z   Pu  s�  I   
I  �*  >�  �;  ��~var ��
  Ec  Cc  	  ��  Oc  Mc  
�  �   val �  [c  Wc  %�  I   �I  ��    ��  #   �	!!  �I  lc  jc  �I  xc  tc   q<  �   �  �	!  <  �c  �c  q<  ��   ��     �<  �c  �c  ñ  �<  Pv Ru    �<  =�   �  ��!  �<  �c  �c  R�  �<  Pv Ru   <<  r�    �  �."  X<  �c  �c  L<  �c  �c  "d<  �  e<  d  d  D  ��   �  �3D  9d  -d  )D  pd  hd     <  �  ��"  0#<  0<  "/<  �  0<  �d  �d  D  ��   �  �3D  �d  �d  )D  �d  �d     D  �  �*�"  3D  e  e  )D  Je  Be   D  ٺ  9   �-�"  3D  oe  ke  )D  �e  �e   q<  �     �E#  <  �e  �e  q<  ��    ��     �<  �e  �e  �  �<  Pv Ru    �<  A�     �#  �<  �e  �e  N�  �<  Pv Ru   J  c�     ��#  "J  �e  �e  J  �e  �e   J  �   �  3   ��#  "J  �e  �e  J  f  f   q<  ��   !  �A$  <  f  f  q<   �    �     �<  .f  ,f  -�  �<  Pv Ru    �<  ջ   ,  �{$  �<  :f  6f  �  �<  Pv Ru   �  ��   7  ��*  �  ]f  If  �  �f  �f  7  �  ng  Rg  �  �g  �g  @�  ��~�  =h  /h  �  uh  sh  �<  ��   j  �'%  �<  �h  }h  �  �<  Pv Ru   D  �   z  �
X%  3D  �h  �h  )D  �h  �h   q<  :�   �  ��%  <  �h  �h  q<  ��   ��     �<  �h  �h  ��  �<  Pv Ru    �<  c�   �  ��%  �<  �h  �h  p�  �<  Pv Ru   D  �  *&  3D  �h  �h  )D  i  i   �<  ��   �   U&  �<  i  i  U�  �<  Pv Ru   D  ��  -   �*�&  3D  &i  "i  )D  <i  :i   D  ��  +   &�&  3D  Hi  Di  )D  `i  \i   q<  �   �  		'  <  ui  qi  q<  ��   ��     �<  �i  �i  ��  �<  Pv Ru    q<  ��   �  o'  <  �i  �i  q<  �   �     �<  �i  �i  )�  �<  Pv Ru    �<  ��   �  �'  �<  �i  �i  ��  �<  Pv Ru   D  V�   V�  :   	�'  3D  �i  �i  )D  j   j   D  �  (	(  3D  Ej  ?j  )D  yj  sj   D  �  	4(  3D  �j  �j  )D  �j  �j   D  �  	_(  3D  �j  �j  )D  �j  �j   D  �  	�(  3D  �j  �j  )D  �j  �j   D    	�(  3D  �j  �j  )D  �j  �j   D    	�(  3D  �j  �j  )D  k  k   D    ")  3D  k  k  )D  k  k   D  ��     	:)  3D  !k  k  )D  +k  )k   :�  $  b)  �  9k  3k  �  Rk  Pk   D  9  +	�)  3D  \k  Zk  )D  fk  dk   D  A�     /	�)  3D  pk  nk  )D  zk  xk   <  �   D  91*  #<  �k  �k  <  �k  �k  "/<  D  0<  �k  �k  D  �    O  �3D  �k  �k  )D  /l  'l     ��  �  E*  Pu  ��  �  ��  �  n�  �  ��  �  ��  c  ��  ;  G�  o  x�  �  ��  �G  ��  D  �*  P��{R��   ��  q  ��  qH  q�  H    B�  I   
�  �+  	�  �  cl  ]l  q<  B�   �  �W+  <  �l  }l  q<  �   �     �<  �l  �l  ��  �<  Pv Ru    �<  p�   �  ��+  �<  �l  �l  N�  �<  Pv Ru   D  ��  :   �.�+  3D  �l  �l  )D  �l  �l   l�  �  Pu   
�  #.  arr �  �l  �l  
�  *-  	�  �  �l  �l  �<  �   �  �E,  �<  m  m  ��  �<  Pv Ru   D  �  ;   �2t,  3D  m  m  )D  1m  /m   q<  J�   �  ��,  <  =m  9m  q<  ��   ��     �<  Nm  Lm  ��  �<  Ps Ru    �<  o�     �-  �<  Zm  Vm  |�  �<  Ps Ru   ۽  �   -  Pu  �  �   q<  ʳ   ʳ     �R-  <  km  im   q<  <�   �  ��-  <  wm  sm  q<  ��   ��  -   �<  �m  �m  ��  �<  Pv Ru    �<  u�   �  ��-  �<  �m  �m  ��  �<  Pv Ru   D  ��      �2.  3D  �m  �m  )D  �m  �m   q�  �E   
  2  obj �  �m  �m  
`  �0  9key �L  ��~
  �.  val �!  n  n  q<  w�   $  ��.  <  *n  &n  q<  g�   g�     �<  ;n  9n  t�  �<  Pv Ru    ��  �  �.  Pu  ��  �   �<  w�   �  �,/  �<  Gn  Cn  ��  �<  Pv Ru   �I  �  �W/  �I  Xn  Vn  �I  fn  `n   q<  ¸   �  ��/  <  �n  �n  q<  �   �  �<  �n  �n  ��  �<  Pv Ru    �<  �   �  ��/  �<  �n  �n  (�  �<  Pv Ru   D  �  �20  3D  �n  �n  )D  �n  �n   D  �  �2A0  3D  �n  �n  )D  o  o   q<  ��     ��0  <  5o  1o  q<  Ծ   Ծ     �<  Fo  Do  �  �<  Pv Ru    �<  ��     ��<  Ro  No  ��  �<  Pv Ru    q<  c�   0  �41  <  co  ao  q<  k�    k�     �<  mo  ko  x�  �<  Pv Ru    q<  ɷ   J  ��1  <  yo  uo  q<  l�   l�     �<  �o  �o  y�  �<  Pv Ru    �<  �   U  ��1  �<  �o  �o  V�  �<  Pv Ru   D  /  �2�1  3D  �o  �o  )D  �o  �o   ��  �F   
�  �2  	  �  �o  �o  b �\   q<  F�   �  ��2  <  �o  �o  q<  �   �     �<  p  �o  )�  �<  Pv Ru    p�    Pu   
h  :3  	  �  p  	p  n �\   q<  ��   }  �3  <   p  p  q<  X�   X�     �<  1p  /p  e�  �<  Pv Ru    ն    03  Pu  �  H   �<  Z�   3  t3  �<  Ap  9p  a�  �<  Pv Ru   q<  ��   >  ��3  <  bp  ^p  q<  ��   ��     �<  sp  qp  �  �<  Pv Ru    q<  D�   d  	04  <  p  {p  q<  R�    R�     �<  �p  �p  _�  �<  Pv Ru    q<  ��   t  	�4  <  �p  �p  q<  ��    ��     �<  �p  �p  ��  �<  Pv Ru    D  p�    p�  6   �4  3D  �p  �p  )D  �p  �p   q<  ��     !5  <  �p  �p  q<  ӹ   ӹ     �<  �p  �p  �  �<  Pv Ru    D  �    �  4   �V5  3D  �p  �p  )D  q  q   D  :  �5  3D  .q  ,q  )D  8q  6q   D  E  �5  3D  Bq  @q  )D  Lq  Jq   D  P  �5  3D  Vq  Tq  )D  `q  ^q   D  [  "6  3D  jq  hq  )D  tq  rq   q<  ɴ   f  #`6  <  �q  |q  q<  �   �     �<  �q  �q  �  �<  Pv Ru    �<  �   q  $�6  �<  �q  �q  �  �<  Pv Ru   q<  ��   �  <�6  <  �q  �q  q<  ��   ��     �<  �q  �q  �  �<  Pv Ru    D  �   �  ;)7  3D  �q  �q  )D  �q  �q   D  �   �  ^Z7  3D  r  r  )D  Gr  Ar   D  ��     }�7  3D  er  _r  )D  �r  �r   q<  ��   -  ~�7  <  �r  �r  q<  u�   u�     �<  �r  �r  ��  �<  Pv Ru    D  G  �8  3D  �r  �r  )D  �r  �r   D  R  �?8  3D  �r  �r  )D  �r  �r   D  ]  �j8  3D  �r  �r  )D  s  �r   D  ��     ��8  3D  s  	s  )D  s  s   q<  ��   �  �8  <  !s  s  q<  ,�   ,�     �<  2s  0s  9�  �<  Pv Ru    q<  �   �  U9  <  >s  :s  q<  ��   ��     �<  Os  Ms  ��  �<  Pv Ru    �<  ��   �  =�9  �<  [s  Ws  Ŀ  �<  Pv Ru   D  �  >.�9  3D  ns  js  )D  �s  �s   q<  ��   �  _:  <  �s  �s  q<  ��   ��     �<  �s  �s  �  �<  Pv Ru    D  �  "*C:  3D  �s  �s  )D  �s  �s   D  �  "Gn:  3D  �s  �s  )D  �s  �s   �<  ��   �  `�:  �<  �s  �s  ��  �<  Pv Ru   D    a.�:  3D  t  t  )D  t  t   ֯  I  �  qH  H�  �  �:  P��|H f�  �G  ��  �H   �   ;  -    !w  �  �;  �  �-�  5	  �A  *op �S�  n   �c  �  ��  l �	\   r �	\   I�;  �  ��;    �  n �\   i �\   neg �\      I�;  lb �\   rb �\    lb �\   rb �\     �  <  F-   � !�  ��  <<  �  �2�  �  �F�  i �\     !#  ��
  q<  �  �2�  �  �F�  i �\     [  ��<  �  �$�   !�  ��  �<  �  �(�   ?@  '�  $�  f  �	D  (�  '$�  Ft  .t  9tok *�  ��}c .
�  �t  �t  
\
  �=  i 9\   �u  �u  num :\   �u  �u  -E  [�   l
  ;L=  <E  v  v   tD  ~�   ~�     ;l=  0�D   	E  ��    |
  =E  v  v  |
  #E  1v  -v     
�
  ?  	m  F�  Jv  @v  i H\   �v  xv  
�
  ~>  ch J�  �v  �v  	E  U�   �
  J">  E  w  	w  �
  #E   w  w    -E  n�    n�     KJ>  <E  1w  /w   	E  �   �
  LE  =w  9w  �
  #E  Pw  Lw     	E  �   �
  F�>  E  cw  _w  �
  #E  zw  rw    -E  #�   �
  I�>  <E  �w  �w   	E  ��   �
  V(E  �w  �w  �
  #E  �w  �w     
�	  J@  i ]\   �w  �w  -E  �   �  	   ^P?  <E  x  x   >D  ��   ��  1   ^�?  ND  x  x  YD  ��   ��  %   �?  iD  x  x   tD  �    �     0�D    �D  *�   �	  c@  �D  .x  $x  "�D  �	  �D  Wx  Ux  "�D   
  �D  dx  `x  �D  yx  sx     \	E  
  _E  �x  �x  
  #E  �x  �x     

  XA  len j\   �x  �x  JÛ    9op l	D  ��}
&
  �@  i m\   �x  �x   J�  �   i p\   )v�  O   �@  j t\   
y  y  	E  |�   A
  t3E  'y  !y  A
  ;#E     D  1
  q$A  3D  Gy  Cy  )D  Zy  Vy   �I  X�   X�     s�I  oy  ky  �I  �y  �y      �D  A�   	  (eC  �D  �y  �y  "�D  	  �D  �y  �y  4-E  T�   +	  ��A  <E  �y  �y   ]	E  @	  ��A  0E  @	  #E  �y  �y    "�D  P	  �D  �y  �y  4	E  �   [	  �)B  E  	z  z  [	  #E  z  z    4	E  /�   f	  �_B  E  3z  /z  f	  #E  Fz  Bz    :�D  v	  	C  �D  az  Wz  4	E  B�   �	  ��B  E  �z  �z  �	  #E  �z  �z    A-E  T�   T�  	   �&�B  <E  �z  �z   K	E  �   �	  �E  �z  �z  �	  #E  �z  �z     4	E  ��   �	  �?C  E  �z  �z  �	  #E  {  {    3-E  ��   ��     �<E  -{  +{      -E  ��   �	  .�C  <E  9{  5{   tD  ��   ��     7	�C  �D  J{  H{   YD  ��   �	  [	�C  iD  X{  R{   	E  ݙ   Q
  |E  s{  o{  Q
  #E  �{  �{     �  D  -    !�  "\   >D  *a "�  *b ".�   !�  \   YD  *c �   !�  \   tD  *c �   !�  \   �D  *c �   !�  \   �D  *str #�  i \   k �  s �     5#  �	E  $�  �&�  +c ��  ^j  ��  +c2 ��      <�  ��  -E  $�  � �  +c �
�   <�  ��  HE  $�  � �   5�  �iE  $�  �!�  $  �4�   L)  �Ħ  #   ��E  �  �!  �  L�  ô�     ��E  �  �  �  ,�  �  T�  ^   ��F  �  �'�  � -val �  �{  �{  )o�  ?   |F  .[  ��F  �N .s  �\   �o 3�I  ��   ��     ��I  �{  �{  �I  �{  �{  �I  �{  �{  �I  �{  �{  8�I  ��     �I  �{  �{     i�  ]I  P�   I  �F  -   ? ,�  �  �  a   �}G  �  �(�  � -val �  B|  >|  )�  B   kG  .�  �}G  �o .;  �\   �� 3�I  9�   9�     ��I  S|  Q|  �I  `|  ^|  �I  m|  i|  �I  �|  |  8�I  9�     �I  �|  �|     �  ]I  P�     �G  -   ? ,�  �  ��  4   �H  �  �(�  � �  �<�  �-val �  �|  �|  A�I  ��    ��     �	H  �I  �|  �|  �I  }  }   ��  ]I  P�   ,�  �  t�     �qH  �  �(�  � �  �4\   �-val �  }  }  }�  ]I  P�   ,_  �  P�  "   ��H  �  �)�  � �  �5\   �-val �  }  }  Y�  ]I  P�   ,Q  �  <�     �I  �  �&�  � -val �  "}   }  E�  ]I  P�   ,�  y  (�     �]I  �  y+�  � -val z  ,}  *}  1�  ]I  P�   <�  k  �I  $�  k-�  +val r   5=  �I  1ptr �  1val &\   1num /\   +p �I  +i \     @   5�  �I  $�    1src /�   <V  \   J  1s "�  +len 	\    5  .J  $�    1src /�   %D  D�  <   �\J  )D  <}  4}  3D  ]}  Q}   %]I  ��  �   �GK  lI  �}  ~}  wI  �}  �}  A�I  ��   ��     s�J  �I  �}  �}  �I  �}  �}  �I  �}  �}  �I  �}  �}  8�I  ��     �I  �}  �}    3]I  �    �  /   klI  ~  ~  ;wI  K�I   �    �  n	�I  /~  +~  �I  E~  C~     %�<  ��  @   �~K  �<  W~  M~  ��  �<  Pv Rw   %q<  ̝  [   ��K  <  �~  ~  q<  �    �     �<  �~  �~  �  �<  Pv Rs    % ;  Ğ  )  �xP  <;  %  �~  H;  ?�  '�  S;  ʁ  ā  _;  �  �  k;  .�  "�  u;  u�  e�  0;  ��  ��  D  �   �  4   �	|L  3D  т  ͂  )D  �  �   :;    �M  @�;  ��{�I  ��    ��     ��L  �I  ��  ��  �I  
�  �   :�;    DM  @�;  ��{�;  /�  #�  �;  p�  ^�  J  >�    >�  %   �,M  "J    ��  J  ΃  ʃ   "�;     �;  �  ��    J  �    �  2   �yM  "J  �  �  J  #�  �   �  �G   D  +  �	�M  3D  6�  2�  )D  I�  E�   D  8�     �	�M  3D  Z�  X�  )D  d�  b�   D  ;  �	N  3D  n�  l�  )D  x�  v�   D  F  �	3N  3D  ��  ��  )D  ��  ��   D  Q  �	^N  3D  ��  ��  )D  ��  ��   D  \  ��N  3D  ��  ��  )D  ��  ��   D  g  �	�N  3D  ��  ��  )D  Ȅ  Ƅ   D  ��    r  �)�N  3D  ڄ  Є  )D  �   �   D  �     �O  3D  �  �  )D  �  �   M�;  ~�  t   AO  ;�;  �;  )�  '�  ޤ  qH   M�;  �  l   nO  ;�;  �;  3�  1�  ]�  qH   u�  H  ��  H  ��  qH  ��  qH  ̣  qH  �  D  �O  P��{R"�   1�  D  �O  P��{R��   H�  D  �O  P��{R��   _�  D  P  P��{R��   x�  D  6P  P��{R��   �  D  UP  P��{R��   �  I  �  D  PsR� #  %�  l�     ��P  &�  � &�  ���  I   %�  ��  !   ��P  &�  � &�  ���  �   %c  Ю     ��P  &r  � &~  ��  �H   _�  ��     �&�  � &�  ��  H    I ~  H}   :;9I8  4 1�B   I   1�B  4 :!;9I  (   	H}  
 !I  4 :!;9I   :!;9I  4 1  4 :!;9I�B  1R�BX!YW    4 :!;9I   :!;9I8  1R�BUX!YW  I  U  'I  1U  '   :;9I  4 1  .:!;9!' !   :!;9I    ! I/  1U   H }  !.:!;9'I !  "4 :!;9I�B  # :!;9I  $1R�BUX!YW  %$ >  &1  ' :!;9I8  (U  ) :!;9I8  *:;9  +4 :!;9I?  ,! I/  -  . 1  /1  0 :!;9I�B  1.1@z  2:;9!	  34 :!;9I  4.1@|  5.?:!;9!'@|  6 :!;9I�B  7 1  8I �~  9. :!;9!' !  :.?:!;9!@|  ;>!!I:!;9!  < :!;9I8  = :!;9!I  >.?:!;9'I@|  ?4 :!;9!	I!  @H }�  A 1R�BUX!YW!  B :!;!�9I  C.:!;9'I@z  D%  E   F$ >  G& I  H '  I&   J   K 'I  L4 :;9I  M:;9  N:;9  O :;9I8  P>I:;9  Q  R 1R�BXYW  SH}�  T.?:;9'   U. ?:;9@|  V.:;9'@z  W.:;9'@|  XH}�  Y1UXYW  Z.1@|  [1XYW    I   :;9I8   !I  H }  'I  '  4 :!;9I�B  4 :!;9I�B  	 :!;9I  
I  ! I/   :!;9I  4 :!;9I�B   :;9I  4 :!;9I�B  $ >  U   1�B   :!;9I�B   :!;9I8   :!;9I   :!;9I�B  U   :!;9I  :;9  4 :!;9I?  4 :!;9I  4 :!;9I     :!;9I�B  :;9!	   .?:!;9!'I@|  !1R�BUX!YW  "  #.?:!;9!'@|  $.?:!;9'I@|  %.?:!;9!'@|  & :!;9!
I8!   '1R�BUX!YW  (.?:!;9!@|  )4 :!;9!	I  * :!;9!I8  +.?:!;9!'@z  ,H}�  -I ~  . :!;9I  /.?:!;9!'@  0.?:!;9'I@z  1 1  24 1�B  34 1  4%  5   6$ >  7& I  8 '  9&   :   ; 'I  < :;9I8  =4 :;9I?<  >4 :;9I  ?4 G:;9  @.?:;9'I@z  A4 :;9I  BH }�  C.?:;9   D.?:;9'@  E. ?:;9@|  F:;9  G :;9I  H.?:;9'@z  I :;9I�B  J.?:;9'   K4 :;9I  L.:;9'I   M :;9I  N.1@z  O1R�BXYW  P.1@|    1�B  I ~  H}  1R�BUX!YW  H }  1UX!YW  4 1�B  1R�BX!YW  	4 :!;9I�B  
U  H}  4 :!;9I�B   :!;9I   :!;9I   :;9I8  I  1R�BX!YW  ! I/  4 :!;9I  (    :;9I8  1R�BUX!YW   :;9I   !I  1X!YW  U   :!;9I8  4 :!;9I     :!;9I  .?:!;9'I@z   $ >  !.:!;9'I !  "1U  # :!;9I  $ :!;9I  %.1@z  & 1  ' :!;9I  ( :!;9I�B  )  * :!;9I  +4 :!;9I  ,.?:!;9!'I@z  -4 :!;9!I�B  .4 :!;9I  /.?:!;9!'@z  0 1  1 :!;9I  2:;9!	  31R�BX!YW  41R�BUX!YW  5.:!;9!' !  6.?:!;9!'I  7.?:!;9!'I !  81  94 :!;9I  :1U  ;4 1  <.:!;9'I !  = I  >4 :!;9I  ?.:!;9'I@z  @4 1  A1R�BX!YW  B>!!I:;9!  C:!;9!  D:!;9!	  E :;9I8  F! I/  G1X!YW!  HH}�  I  J  K1R�BUX!YW  L.?:!;9!'@z  M1  N%  O$ >  P:;9  Q:;9  R& I  S'I  T:;9  U   V'  W 1  X 1  YI �~  Z.:;9'I@|  [.:;9'   \1UXYW  ]1UXYW  ^4 :;9I  _.1@z   �E            ����P����U  ����0�����1�����2�����3�����4�����5�����6�����7�����8�    ����0�����0�   ����V    ����x�����x�     ����P����P   ����P        ����D�����D�����D�����D�                             ����W����	��  4$�����W����	��  4$�����W����W����	��  4$�����W����	��  4$�����W����	��  4$�����W����	��  4$�����W����	��  4$�        ����:�����:�����:�����:�            ����0�����S����S����S����S����S            ����s 
�� "�����s
�� "�����s 
�� "�����s 
�� "�����s 
�� "�����s 
�� "�           ����P����	rw #D�����
r�}w #D�����r�}��  4$#D�����	rw #D�                ����s 
�� "#
�����s
�� "#
�����s 
�� "#
�����s 
�� "#
�����s 
�� "#
�����s 
�� "#
�����s 
�� "#
�����s 
�� "#
�        ����@� �����@� �����@� �����@� �        ����
 �����
 �����
 �����
 �                   ������{�����V������{�����V������{�����V������{�����V������{�           ����P������{������{������{������{     ����@� �����R  ����	r ?� �����r ?� �-( �     ����P����W   ����P     ����@� �����@� �����@� �����@� �����@� �     ����
 �����
 �����
 �����
 �����
 �         ������}�����W������}�������}�������}�����W������}�       ����R����V����R  ����V  ����	v @� �����v @� �-( �     ����P����p�����P       ����P����P����U   ����P  ����	p ?� �      ����
 �����
 �����
 �      ����W����W����W        ����V����V������{�������{�         ������{�����Q����U����U                    ����0�����R����v�����V����v�����R����v�����R����v�����V����v�      ����0�����R����R        ����0�����Q����12q 0)( �����12q 0)( �����Q    �B�PL��P�XL�    �C�Px��P�Xx�        �C�C� �C�ES�O�OS�X�X�       �E�Ou#��O�Pu#��P�Xu#�         �J�KW�K�Ou#D��O�Pu#D��Q�Xu#D�         �J�JP�J�Ou�}�O�Pu�}�Q�Xu�}         �J�KS�K�Ou�}�O�Pu�}�Q�Xu�}      �K�O@��O�P@��Q�X@�         �K�KP�K�Ou�}�O�Pu�}�Q�Xu�}       �C�C0��E�Ew��E�EW�X�X0�     �D�DP�D�Eu�}�O�Ou�}       �D�DR�D�Eu�}�O�Ou�}  �I�Ip� 3$u�}"�            �K�K0��K�Ku�}�L�LP�L�Ou�}�Q�QP�V�Xu�}      �K�Ku�}4�I "��L�Ou�}4�I "��V�Xu�}4�I "�     �L�NW�V�XW  �V�Vu�}4�I "      �V�VP�V�VQ�V�Xu�}  �V�Wu�}  �V�Vu�}4�I "  �V�XW  �M�Nu�}4�I "     �M�Ms�M�Ou�}   �M�Ms     �M�NP�N�Ou�}     �M�Ms�M�Nu�}     �M�NR�N�Ou�}   �M�NW    �M�NP�N�Ou�}               �O�OQ�O�Pu�}�Q�Q0��Q�Tu�}�T�TQ�T�Vu�}�X�Xu�}      �Q�Tu�}
��} "��T�Vu�}
��} "��X�Xu�}
��} "�         �O�OS�Q�TS�T�VS�X�XS                  �Q�Ru�}w�D��T�U
u�}p D��U�Uu�}w�D��U�Uu�}w�D��U�U
u�}p D��U�Vu�}w�D��X�Xu�}w�D��X�X
u�}p D��X�Xu�}w�D�                 �Q�RR�R�Tu�}�U�Uu�}�U�UR�U�Uu�}�V�VP�X�Xu�}�X�XP           �R�RR�R�Tu�}�U�Uu�}�U�UR�X�XR          �R�Rp 8��R�Tu�}�U�Uu�}�U�Up 8��X�Xp 8�    �R�RP�U�UP         �S�Sp 3$��S�SP�S�St �S�Su�}         �O�PP�P�PQ�X�XP�X�XQ        �P�P��  p q @��P�P��  u�}q @��X�X��  u�}p @��X�X��  u�}q @�        �P�Pp q ��P�Pp q D+( ��P�Pu�}q D+( ��X�Xu�}p D+( ��X�Xu�}q D+( �       ����U����U�����    ����P       ����Q����
@�  r "�����	r @� �����	r A� �     ����P����R  ����W       ����P����R�����\         ����P����R����	p @� �����
@�  p "�����	p @� �           ���0�����0�����W����w�~�����0�      ��ųPų̳��  ����P  ����   ����0� ���0�  ����5 �            ͳڿ
�����
�����
�����
�����
�����
�            ͳڿ
������
������
������
������
������
��                                              �ݴ0�ݴϿ��}������}������}������}����V����Q������}����Q������}������}����Q������}����R������}����Q����P������}����V������}����V������}������}                                          �ݴ0�ݴƺ��}ƺɺPɺ���}����}�����}������}��Ͽ��}������}����P������}������}����P������}����P������}������}������}������}������}������}������}������}������}����
s�	��}"�����P����
s�	��}"�����V������}����
s�	��}"�                      �ݴ@�ݴ����}��̵Q̵����}����Q��Ͽ��}������}������}������}������}������}                  �ݴ0�ݴϿ��}������}������}������}������}������}������}������}                          �ݴ0�ݴ����}ֻϿ��}������}������}������}������}������}������}������}������}������}������}            �ڿ
������
������
������
������
������
��                            �ݴ0�ݴ����}ֻϿ��}������}����P������}������}������}������}������}������}����Q������}������}                            �ݴ0�ݴ����}ֻϿ��}������}����P������}������}������}������}������}������}����R������}������} 	                                   �ݴ0�ݴϿ��}������}����0�������}������}������}����0�����P������}������}����0�����P������}����0�������}������}����0�������}                  �ݴ0�ݴϿ��}������}������}������}������}����P������}������}                                 ����S����P����S������}��ֻSֻ���}���S��Ͽ��}ϿڿS����S������}����S����S������}����S����S               ����P������}ֻ���}��Ͽ��}����P������}������}             ����P������}ֻ���}��Ͽ��}������}������}             ����0�����VͺպSٺ�Vֻ�S��ϿV����0�             ����0�����Wͺպ0�ٺ�Wֻ�0���ϿW����0�      ��
v 2#p ����
v 2#r �����
v 2#r �                     ����0�����R����s���ζSζ�R�ٺs�ٺ�Sֻ�s�����R��Ͽs�����s�����s�       ����r 
��} "���ĸ��}
��} "�������}
��} "�     ������}������}     ���W����W     ����p 
�� "������� 1
�� "� ̵�V ̵���}  ��P                 ����P��μs�	����s�	����s�	����s�	����s�	����s�	����s�	     ���q 
��} "�������}
��} "�  ��ѽP   ̽����}                 ����P����s�	����P����s�	����P����s�	����s�	����P                 ����Q����s�	����Q����s�	����Q����s�	����Q����s�	      ����0�����P����P����P  ������}  ����
��  ����0�   ����s�	     ����R����R   ����Q     ����p 
��} "������} 1
��} "�     ����p 
��} "������} 1
��} "�     ����p 
��} "������} 1
��} "�       ����q 
��} "������} 1
��} "�����q 
��} "�       ����	v w q "�����P������|     ��� �  ����� �  ����� �  �     �����  �������  �������  �      ���W����W����W      ���� ����� �����           ���	������S����S����S����R          ���	������V����V����V����V  ����s 
�@% "�        ���0�����R����R����R    ����W����w�~�                   �"�"P�"�$S�$�$�\p "2$p "2$�I "�$�%�\`I "2$`I "2$�I "�%�%
�� &�-� ��%�%S�%�%�\p "2$p "2$�I "�%�%�\p "2$p "2$�I "�%�%S                   �"�#R�#�$w �$�$�\p "2$p "2$�I "�$�%�\`I "2$`I "2$�I "�%�%
��&�-� ��%�%�\p "2$p "2$�I "�%�%�\p "2$p "2$�I "�%�%�\p "2$p "2$�I "�%�%w                    �"�#Q�#�$w�$�$�\p "2$p "2$�I "�$�%�\`I "2$`I "2$�I "�%�%
��&�-� ��%�%�\p "2$p "2$�I "�%�%�\p "2$p "2$�I "�%�%�\p "2$p "2$�I "�%�%w      �#�$p 4�I "��$�%`I 4�I "��%�%p 4�I "�               ܝ��P��ɟSɟͧ
�� &�-� �ͧ��S��ݨ
�� &�-� �ݨ�S���
�� &�-� �               ܝ��R��ʠUʠͧ
��&�-� �ͧ��U��ݨ
��&�-� �ݨ��U����
��&�-� �               ܝ��Q��ʠ��{ʠͧ
��&�-� �ͧ����{��ݨ
��&�-� �ݨ����{����
��&�-� �           ����P����R������{ͧԧPݨ�P���R            ����P������{��ͧ��{������{��ݨ��{������{                            �ΠUΠ�S���U����S����U��֤u�֤�R�ĦUĦǦu�ǦզQզ��U��ͧU����U��ȨU����U              ����u s �����P������{����u s �����P������{Ħ����{������{       Ǧ�P���q����q    Ǧ��Q����Q          ��u q ����P������{����P����r�      ����u r �����P������{  ����	s  : "�  ����V ����1�    ����P������{    �����{Ȩݨ��{    ���d� Ȩݨd�      �����{Ȩݨ��{     ���d� Ȩݨd�                                                                                                                                                d�R��P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��	
��&�-� ��	�
P�
�
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P��
��&�-� ���P�� 
��&�-� �� � P� �!
��&�-� ��!�!P�!�"
��&�-� �         d�Q��
��&�-� ���Q��"
��&�-� �         dzp z�u ��p ��"u           PGWHSWTcW                2R2;Q;BRHTRTXQX\r�\cR     5PHPP     *2QHTQ                     �%�%P�%�%S�%�%s��%�&S�'�-S�-�-S�-�-V�-�-Q�-�.vx��.�.vx��/�1S         �&�'R�.�/R�/�/R�/�/R         �&�&0��&�&P�&�&P�/�/0�       �&�&0��&�&Q�'�'Q       �.�.0��.�.V�.�/V       �-�-P�-�.W�.�.W      �-�-0��-�.P�.�.P        �-�-0��-�-vw q "��-�.q v #	��.�.vw q "��.�.q v #	��.�.vw q "�                 �-�-R�-�-r0��-�.q �.�.q�.�.R�.�.r� ��.�.R�.�.r7�     �1�1P�1�2Q         �1�20��2�2P�2�2P�2�2P         �2�2P�2�2
�� &�-� ��2�2P�2�2
�� &�-� �             �2�3P�3�3S�3�3
�� &�-� ��3�4S�4�4
�� &�-� ��4�4S     �3�4S�4�4S                 �4�5P�5�5S�5�5
�� &�-� ��5�>S�>�>
�� &�-� ��>�>S�>�>
�� &�-� ��>�BS     �5�>S�>�BS       �X�YP�Y�Y�P�Y�ZQ�Z�\�P               �X�YR�Y�[U�[�\
��&�-� ��\�\R�\�\U�\�\
��&�-� ��\�\U         �Y�YR�Y�[U�[�\
��&�-� ��\�\U       �Y�Y�P�Y�ZQ�Z�\�P�\�\�P     �Y�\1��\�\1�      �Z�ZP�Z�\�T�\�\�T   �Y�Y0� �Y�Z2�    �Z�ZP�Z�Z�T  �[�[�T�\�\�T  �[�[R�\�\R  �[�[�T�\�\�T  �[�[R�\�\R   �[�\U       �\�\P�\�\S�\��
�� &�-� �     �\�\R�\����}       �\�\P�\�^S�^��S     �]�]R�^�^R         �]�]0��]�^R�^�^R�_�_0�      �^�^��~��^�^P�^�^��~�      �^�_��~��_�_P�_�_��~�      �_�`��~��`�`P�`�`��~�  �c�cW  �d�dW  �e�eW      �f�f��~��f�fP�f�f��~�      �g�g��~��g�gP�g�g��~�      �g�g��~��g�gP�g�g��~�      �g�h��~��h�hP�h�h��~�      �h�h��~��h�hP�h�h��~�      �h�i��~��i�iP�i�i��~�                �i�i0��i�jR�j�jr��j�jR�j�j��}�k�kR�o�oR�o�oR          �i�i��~��i�jW�k�kW�o�oW�o�oW        �j�j��~��j�jP�j�j��~��j�j��~�           �p�pW�q�qW�r�rW�r�sW�s�sW  �s�sW      �k�k��~��k�kP�k�k��~�        �l�l0��l�l��}�l�mQ�m�o��}          �l�l��~��l�mW�m�mW�n�nW�n�nW  �m�mW      �o�p��~��p�pP�p�p��~�      �p�q��~��q�qP�q�q��~�      �q�q��~��q�qP�q�q��~�      �r�r��~��r�rP�r�r��~�      �t�t��~��t�tW�u�uW      �v�v��~��v�wW��ЅW      �w�w��~��w�wP�w�w��~�      �w�x��~��x�xW����W          �x�y��~��y�zW���W����W��W      �z�z��~��z�{WЅ�W      �{�{��~��{�}W��րW    �}�}��~��}�~W      �~�~��~��~�~P�~�~��~�      �~�~��~��~�~P�~�~��~�  ��W         ����WӃ�W����W��҄W      ������~�����P������~�      Ӂ���~���P����~�      ������~�����P������~�      ��ʂ��~�ʂ΂P΂ς��~�      �����~�����P������~�               ����W��ӃW���W����Wڄ�W����W���W  ����W                             ؆�R���P����R����V��ʇ��Wʇ�S���s�����S��ی��Wی�R�����W����s�������W��Ώs�Ώ����W             ��ʇPʇ܇U܇�P���U����U��ΏU                ��ʇ0�ʇ͇q�͇Їq�Ї�Q���q�����Q����q���Ώq�              ������_�����U��ی��_�����_�������_�������_�Ώ����_�     ̈P̈��V                                                  ���U������W������W#�����V��ω��WωیS����W����S������W������W#�������W��ɍRɍލ��Wލ��S������W����S������W����Q��Ďq�ĎҎQҎ����WΏڏSڏ����W���S�����W������W#�������W#�����V����R����S������W    ����0�����0�����1�           Ǎލ0�ލ�R���0�Ώ��R����R       ����0���ҎS����0�ڏ�0�����0�           ����P����Q������W������Wؙ����W        ����R������W������Wؙ����W ����1�    ���P������W                          ݑ����[�����Q����V����S����V����S��͖V͖�v���V���W���Vؙۙv�ۙ�Q���V            Ғ֒v s �֒�P����W����v s ���ɖPɖ����Wؙ����W        ����w v �����P������W����w v �     ۙ��P����q  ۙ��Q      ���v q �����P������W  ӛ��	s  : "�  ӛ��U     ��ȕ��W�����W     ��ȕP���P     ��ȕ��W�����W     ��ȕP���P     ����P����P           ��V���v���׋V׋܋q,܋ʌ��W#,������W#,    �یU����U ���2�  Ҋ�U ����U ����P    ��یU����U        ��ҌPҌیd� ����P����d�                      ����P���V��
�� &�-� ����V����
�� &�-� �����V����
�� &�-� �����V����
�� &�-� ���ٝV       ��МP���P����P       Ĝ�V����V����
�� &�-� �     ʜ�S����S              ߪ��0���ҫWݫ�W���w�����W����1�����W��ήWή׮0�׮°W            ߪ��0���ҫ��[ݫ����[����0������[��q����Q��°��[            ߪ��0�����U����0���ҫUݫ��U����u�����U��°U              ߪ����  ���ҫVݫ��V����V����v�����V����v�����V����v���°V                                                  ����P��ūPݫ��P����	� w "
`����	� w "
a����P����P������[����P����	� u "
 ��ƭ	� u "
!ƭ�P��	� q "
 ���� ��["
 ����	� q "
!����P����P��ЮP׮�P���P��ůP��P����P����P����P    ����@� �����@� �           ����0�����
@�  p "�����
@�  p "�����	p @� �����	p A� �����
@�  p "�               ����0�����U����U����U����U����u�����V����U        ����R����R����R����R    ������}�����Q    ������{�����P    ����@� �����V    ����W����P       ����P����� �����        ����0�����V����v�~�    ����V����v�~� �
            �/�/P�0�0P                   �+�,P�,�,
� 
�1&��,�,P�,�-
� 
�1&��-�.P�.�.p�}��.�.
� 
�1&��.�.P�.�.
� 
�1&�        �+�+
�
,1&��+�+w 1&��+�,
�
,1&��,�.
�
,1&�    �,�-�
,1&#(��.�.�
,1&#(�      �,�,ȟ�,�,V�.�.ȟ   �-�.V    �,�-	�u D��.�.	�u D�         �,�,
r �2 "��,�-R�-�-�2 �.�.R    �+�+� 
���+�+P �+�+�
,�             �"�"Q�"�#�H�#�%�D� "��%�*�
�1&� "��*�*�D� "��*�*�
�1&� "�         �"�"R�"�$�T�$�*�
,1&�"��*�*�
,1&�"�         �$�&V�&�*�T#(��*�*V�*�*�T#(�    �$�%ȟ�*�*ȟ    �%�*D��*�*D�         �'�(Q�(�)�L�)�*�T#���*�*�T#��        �%�&0��&�&�D�&�&P�&�(�D     �&�&V�&�(V            �&�&w~��&�&wj��'�'w~��'�'P�'�'���'�'w~�   �&�&Q �!�!�
�� �"�"�
,�         ��P��W�!�!P�!�!W   ��P     ��� ���      ������    ��@���@�         ��P��V���X���X��V             ��P��R���L���L��P��R          ��0����D��R���D��0�       ��w 1���W��W    ��0���0�     ��P���\   ��P   ��Q     ��� ���            �����S�����S���       �����R��R     �����Q     ��� ���            �����S�����S���       �����R��R     �����Q    ��0���S        ��S��S������S           ��U��P��U���\��U       ��P��V��V       ��S��	DJ 1���S      ��0���P��0�     ��P���@     ��V�	�	V         ��	V�	�	v{��	�	P�	�V     ��	U�	�U          �	�	P�
�
P�
�
p��
�
q��
�
q p "#��
�q p "#�        �
�
P�
�
p��
�
q��
�
q p "#��
�
q p "#�    �
�
0��
�P    �
�
0��
�
P   ���     ��P��P   ��P     ��P��V   ��P  ��p v ���p v O-( �   ��P       ��V��P��V     ��P��R       ��p v ���r v ���u�v �-( ���r v �-( �           ��� ��Q��� ��Q���            �����V�����V���           �����S�����S���      ��0���P��P    ��0���U       ��� ��� ���      ��� ��P     �����Q     ozPz�W     ��P��U    ��0���V  5�   5�      0�p � �	p � #�*p � �      ��p 0r 8$"|J "���p 0� 8$"|J "����0� 8$"|J "�   ��R���  ��e�           ��P��p���P��P��P��R��P �4            ����P�����h     ����P�����h     Ą΄P΄Ԅ�h     �0�0� �1�2�           �0�00��0�0W�1�1W�1�1W�1�20�         �0�0R�0�0Q�0�0R�1�1Q      �0�0S�1�1S�1�1S     �1�1��1�1S   �1�1Q   �/�0V      �/�/��/�/��0�0�      �/�/� �/�/� �0�0�         �/�/0��/�/W�/�/W�0�0W         �/�/Q�/�/R�/�/Q�/�/R        �/�/V�/�/S�/�/S�0�0V     �.�/� �/�/S       �.�/��/�/P�/�/�   �.�/v 
P� "#���     �.�.��.�.P   �.�.R       ��łPłւS���P  ���R  �����y�      ����R����r�����r p "#�����r p "�����r p "#�    ����0�����P  ււ��w������w  �-�.�   �-�.�       �-�.0��.�.p � ��.�.	p � #��.�.	p � #��.�.p � �      �-�-P�-�-P�-�-�#  �,�-P         �+�+0��+�,W�,�,W�,�,W         �+�,R�,�,Q�,�,R�,�,Q      �+�,S�,�,S�,�,S           �)�)0��)�*W�*�+W�+�+W�+�+0�         �*�*R�*�*Q�*�*R�*�*Q      �)�*S�*�*S�+�+S     �*�*��*�*S   �*�*Q      �'�'0��'�'U�'�(0�       �'�'R�'�'R�'�(V    �'�'0��'�'0��'�(1�             �$�$P�%�%P�%�%Q�%�%r 3%��%�&Q�&�&P        �$�$N��$�$M��%�%N��%�&V�&�&��2��&�&N�      �%�%p 0-���%�&�#0-���&�&p 0-��         �{�{P�{�|U�|�|
�� &�-� ��|��U        �{�{P�{�|U�|�|
�� &�-� ��|��U          �{�|u��|�u���u���Ӏu����u�         �|�|P��P�����}Ӏ���}             �}�}P�}�}��}�}�}P�}�}��}���P������}    �|�}U��ӀU   ��΀U   �}�}U���U    �}�~��  ��~�~Q  �~�~S  �}�}U   �~�~��  ��~�~Q   �~�~��}�~�~S    �~�U����U   ����U     �{�{P�{�{U��U  �|�|U��U    �|�|��  ��|�|Q      �|�|P�|�|��}�|�|V    ����  ����S  ���Q    ����UӀ�U   Ӏ�U         �p�qP�q�tU�t�t
�� &�-� ��t�{U      �q�tU�t�t
�� &�-� ��t�{U                 �q�qP�q�t��}�t�tP�t�t��}�t�z��}�z�{��}�{�{P�{�{��}            �q�tu��t�yu��y�yP�y�zp|��z�{u��{�{u�         �q�qP�q�t��}�t�{��}�{�{��}    �t�tU�{�{U   �{�{U     �s�tP�t�t��}    �s�sU�z�{U   �z�zU    �t�tU�z�zU       �y�yP�y�zV�{�{V     �z�zP�{�{P   �{�{R   �q�q��  ��q�qQ     �q�qP�q�q��}�q�qW    �r�rQ�t�tQ    �r�rW�t�tW  �r�rQ  �r�rW  �r�rQ  �r�rW  �s�sQ  �s�sW  �s�sQ  �s�sW  �u�uQ  �u�uW  �u�uQ  �u�uW  �u�uQ  �u�uW  �v�vQ  �v�vW  �v�vQ  �v�vW  �v�vQ  �v�vW  �v�wQ  �v�wW  �w�wQ  �w�wW  �w�wQ  �w�wW  �w�xQ  �w�xW  �x�xQ  �x�xW  �x�xQ  �x�xW  �x�xQ  �x�xW  �y�yQ  �y�yW   �y�yP   �y�yV   �q�qU�{�{U                                                             �3�4P�4�5U�5�5
�� &�-� ��5�6U�6�7��{�7�8
�� &�-� ��8�8P�8�9U�9�9��{�9�:
�� &�-� ��:�;U�;�;
�� &�-� ��;�AU�A�A��|H��A�CU�C�C
�� &�-� ��C�DU�D�D
�� &�-� ��D�D��{�D�SU�S�S
�� &�-� ��S�dU�d�d
�� &�-� ��d�gU�g�gP�g�g��|H��g�iU�i�iP�i�oU�o�p
�� &�-� ��p�pU�p�p
�� &�-� �                                                            �4�4P�4�5U�5�5
�� &�-� ��5�6U�6�7��{�7�8
�� &�-� ��8�8P�8�9U�9�9��{�9�:
�� &�-� ��:�;U�;�;
�� &�-� ��;�AU�A�A��|H��A�CU�C�C
�� &�-� ��C�DU�D�D
�� &�-� ��D�D��{�D�SU�S�S
�� &�-� ��S�dU�d�d
�� &�-� ��d�gU�g�gP�g�g��|H��g�iU�i�iP�i�oU�o�p
�� &�-� ��p�pU�p�p
�� &�-� �                                                                            �4�4P�4�5��{�5�6��{�8�8P�8�9��{�:�<��{�<�=u��=�?��{�A�C��{�C�D��{�D�E��{�F�Fu��G�Gu��G�H��{�I�I��{�I�Iu��J�N��{�O�Ou��O�P��{�Q�R��{�R�S��{�S�S��{�S�T��{�U�[��{�[�\��{�]�]��{�]�_��{�_�`u��`�b��{�d�f��{�f�f��{�f�fP�g�gP�g�gp|��g�gP�g�hp|��j�j��{�j�ju��j�k��{�l�l��{�l�lu��m�mu��n�n��{             �_�_P�_�`��|�`�`P�`�`��|�j�j��|�j�jP   �`�`p Hr "#���     �`�`��{�`�`W   �`�`S       �^�_u��_�_Q�j�ku�           �^�_��~��_�_W�_�_R�j�k��~��k�kP    �_�_U�`�aU   �`�aU   �_�_U�`�`U    �j�j��  ��j�jR      �j�ju��j�js��j�jS         �f�fP�f�gV�g�hV�i�jV           �g�gP�g�g��|�i�i��|�i�iP�i�j��|   �g�g0�     �l�lP�l�m��{     �l�lP�l�lP  �l�m
��      �l�l0��l�l	
���|��l�l	
���|��l�m	
���|�       �l�lS�m�mP�m�mS    �m�m�  ��m�mR    �m�mu��m�mV   �l�lU�m�mU   �9�9V   �9�9V     �9�:P�:�:W   �5�5Q     �5�5��~��5�5P    �5�5U�8�9U   �8�9U  �5�6U�9�9U       �6�7��{�9�9��{�D�D��{         �6�6P�6�7��{�9�9��{�D�D��{        �6�60��6�7W�9�9W�D�DW            �6�6��{�6�6Q�6�6R�6�6Q�9�9R�D�D��{        �6�6V�6�6S�9�9S�D�DV         �7�70��7�7W�9�9W�S�SW            �7�7��{�7�7R�7�7Q�7�7R�9�9Q�S�S��{        �7�7V�7�7S�9�9S�S�SV        �J�J�  ��J�KS�U�US�a�a�  �        �J�J��|�J�KV�U�UV�a�a��|    �K�K6�  ��K�KQ  �K�KV    �K�KU�M�MU   �M�MU  �K�LU�M�MU   �L�L6�  ��L�L7�  �     �L�L��{�L�LP�L�Lp�   �L�LQ    �L�L��{�L�LP    �L�MU�M�MU   �M�MU   �M�MU�M�MU                    �U�Y��{�^�^��{�a�a��{�a�d��{�e�f��{�h�i��{�j�j��{�k�l��{�m�n��{�n�p��{                        �U�YU�^�^U�a�aU�a�dU�d�d
�� &�-� ��e�fU�h�iU�j�jU�k�lU�m�nU�n�oU�o�p
�� &�-� ��p�pU�p�p
�� &�-� �                        �U�YU�^�^U�a�aU�a�dU�d�d
�� &�-� ��e�fU�h�iU�j�jU�k�lU�m�nU�n�oU�o�p
�� &�-� ��p�pU�p�p
�� &�-� �            �V�Y��{�^�^��{�a�au��a�b��{�e�f��{�k�k��{             �V�V0��V�YS�^�^@��a�a0��e�fS�k�k@��k�kS   �p�pU   �U�UU�a�aU   �U�UR�a�a�  �   �U�UQ�a�a��|    �U�VU�a�aU   �a�aU   �V�VU�a�aU    �X�X�  ��X�XQ  �X�XV   �V�VU�X�XU    �V�W�  ��W�WQ  �W�WV    �W�W�  ��W�WR    �W�W��|�W�WV    �W�XU�k�kU   �k�kU    �X�YU�e�eU   �e�eU   �Y�YU�e�fU      �^�^��  ��^�^	v ��  "��^�^	v ��  "��^�^	v ��  "�      �^�^��{�^�^	� v "���^�^	� v "���^�^	� v "��     �a�a	v ��  "��a�b	v ��  "��b�b	v ��  "�     �a�a	� v "���a�b	� v "���b�b	� v "��  �b�bR  �b�bW  �b�cR  �b�cW  �c�cV  �c�cW  �c�cV  �c�cW  �c�dV  �c�dW  �d�dV  �d�dW   �i�iR   �i�iV      �j�j0��j�jR�j�jR   �j�jP  �k�kV  �k�kQ  �m�nV  �m�nQ    �o�p��{�p�p��{      �o�oP�o�p�� &�-� #��p�p�� &�-� #�      �o�o0��o�pW�p�pW        �o�o��{�o�o	� s "���o�o	� s "���o�p	� s "��        �o�oQ�o�oq s "��o�oq s "1��o�pq s "�       �<�<P�<�=��|�S�T��|    �;�<U�I�IU   �I�IU   �<�<U�S�TU    �<�<�  ��<�<Q    �<�<��{�<�<S       �P�PP�P�S��|�Z�[��|   �Q�QP   �Q�QU�R�RU    �Q�Q�  ��Q�QS  �Q�QV    �R�RU�R�SU   �R�SU   �R�RU�S�SU  �=�=U    �O�PU�[�[U   �[�[U    �P�PU�Z�[U    �P�P��  ��P�QQ  �P�QS                 �E�EP�E�I��|�I�J��|�N�O��|�S�S��|�T�T��|�[�[��|�\�\��|   �N�NP    �N�NU�T�TU   �T�TU �F�FU�G�GU   �F�FQ       �F�F��|�F�FR�T�T��|    �F�GU�O�OU   �O�OU    �G�GU�J�JU�N�OU�O�OU    �H�H�  ��H�HQ  �H�HV        �I�I��  ��I�JV�N�NV�O�O��  �      �I�I��{�I�JW�N�NW    �H�HU�S�SU   �S�SU   �H�IU�S�SU  �J�JU   �J�JU    �E�EU�\�\U   �\�\U    �E�EU�\�\U      �E�F��  ��F�FQ�J�JQ    �F�FV�J�JV     �Z�ZP�]�]P    �Z�ZU�]�]U   �]�]U     �C�CP�j�jP    �B�CU�f�fU   �f�fU        �4�4P�4�4U�8�8P�8�8U    �4�5U�=�=U   �=�=U    �C�CU�M�NU   �N�NU  �8�8U   �8�8U    �:�:��  ��:�:Q    �:�:u��:�:V    �:�;U�I�IU   �I�IU    �;�;�  ��;�;Q      �;�;W�;�;��{�;�;V  �=�=Q  �=�=V  �>�>Q  �>�>V  �>�>Q  �>�>V  �>�>Q  �>�>V    �?�?U�S�SU   �S�SU  �?�?U�S�SU    �T�TU�[�[U   �[�[U     �?�?�  ��?�@Q�T�TQ     �?�?u��?�@V�T�TV         �@�@��{�@�@P�@�@��{�U�U�  ��\�\��{     �@�@V�U�Uu��\�\V    �@�@R�]�]�  ��n�n�  �     �@�@v��@�@V�]�]u��n�nu�    �@�AU�f�fU   �f�fU  �A�AQ  �A�AV  �A�AQ  �A�AV  �B�BQ  �B�BV  �B�BR  �B�BV    �D�DU�[�\U   �[�\U    �O�OU�Z�ZU   �Z�ZU  �T�UU�[�[U    �e�e�  ��e�eR    �e�eu��e�eS    �\�\U�]�]U   �]�]U  �Y�YQ  �Y�YV    �Y�ZR�f�fR    �Y�ZV�f�fV  �\�]U�]�]U    �d�d�  ��d�eR    �d�du��d�eV                         ��R��
��&�-� ���R��	��}�	�	
��&�-� ��	�	R�	�

��&�-� ��
�R����}��R����}��R                                         ��P��u ��}"����}��P��w ��	
��}��}"�	�	��}�	�
��}�
�
P�
�
w �
���}��P����}��q0�����}��
��}��}"����}��
��}��}"����}����}        �
�
0��
�S��S��S            �
�
0��
�
V�
�V���`��V��V  �
�
R�
�
R     �
�
R��R     �
�
Q��Q           ����}����}����}����}����}            ��0���W��W��0���W��W                ��P��\���:���P��\���P��P��P��:�    ��R��R     ��P��P   ��R    ��R��R     ��P��P    ��R��R         ��P����}��P����}     ��R��R��R��R    ��R��R     ��r v "��r v "    ��0���s�  ��R   ��V  ��V          ����}���W��Q��W�	�
W  ��0�     ��P�	�
P       ��W��Q�	�
Q     �	�	R��R     �	�	Q��Q            ��	Q�	�	q��	�	Q��Q����}��Q    ��0���P      ��0���Q��Q     ����}����}����}    ��P��P     ����}��W    ����}��S    ����}���Q      ��R��R��R   ��S   ��R��R       ����}��s ����}     ��S��S    ��R��R     ����}��s    ��R��R     ��w ��w            ��Q��Q��:���Q��Q        ��R��R��R��R��R     ��Q��Q  ��R    ��R��R     ��s ��s    ��R��R     ��u p "1��u p "1 ��R  ��R��R ��P      ��P��P��w     �	�	��}����}     �	�	P��P     �"�"P�"�"R  �"�"��  �"�"0�    �"�"P�"�"q�~�    �"�"P�"�"q�~�      �"�"0��"�"	p q #���"�"	p q #���"�"	p q #���"�"	p q #��     �!�!P�!�"R  �!�"
H�  �!�"0�    �!�!P�!�"q�w�    �!�!P�!�"q�w�      �!�!0��!�!	p q #���!�"	p q #���"�"	p q #���"�"	p q #��   ��P     �����S   ��R   ��P   ��P   ��P   ��P          P$P+1P8<P              RS+R+/S/8r�8<R           <\P\�R��P��r�t���
�� &�-� �     p�V��P  p�
�  p�0�  p�V    p�V��P  px0�      ��P��r�t���
�� &�-� �     ����  ���P   ��R           ��P��W��pl���W��pl�           ��P��S��
�� &�-� ���S��
�� &�-� �   ��S                                                                                           ��R��S��
��&�-� ���R��S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��
��&�-� ���S��w|���
��&�-� ���S��
��&�-� ���S��
��&�-� ��� S� � 
��&�-� �� � S� � 
��&�-� �� � S� � 
��&�-� �� � S� � 
��&�-� �� � S� � 
��&�-� �� � S� �!
��&�-� ��!�!S                         ��Q����{��Q����{��
��&�-� �����{��
��&�-� �����{��
��&�-� �����{��
��&�-� ���!��{       ��� ��� ��!�             ��P����{��P����{����{��!��{             ����{����{����{����{����{��!��{                 ����{����{����{����{����{����{����{��!��{   ��!�0;  �   ����  ���W   ����{��U   ��R       ����{���W��P             ��P��P��S��r 3%���S��S            ��?���>���=���>���W��U����{1���U����{2�   ��R     ����{���P      ��p 0-����
��{0-����
��{0-��   ��Q     ��W��P    ��W��W    ��U��U  ��W  ��U  ��W  ��U  ��W  ��U  ��W  ��U  ��W  ��U  ��U  ��W           ��Q��R��Q��R��q�    ��W��W  ��P  ��W   ��U   � � W                  /}              �d       0}                O~       D�  [B                  2HP �&�'�.�.�.�/�/�/ �-�.�.�. �-�-�-�.�.�. �-�-�.�.�.�. �3�4�4�4 �5�>�>�B �C�C�C�C�C�E�O�O �C�C�C�E�O�O�O�O �K�O�Q�Q�V�X �K�K�L�O�V�X �L�L�V�X �O�P�X�X �P�P�X�X �Q�V�X�X �Q�T�T�V�X�X �Y�\�\�\ �[�[�[�[�\�\ �\�\�]�^�^�� �^�^�`�a �^�_�a�a �i�j�k�k�o�o�o�o �j�j�j�j �j�j�p�p�q�q�r�r�r�s�s�s �k�m�m�o �t�t�u�u �v�w��Ѕ �w�x���� �x�z��������� �z�{Ѕ� �{�}��ր ������Ӄ�������ڄ ������Ӄ�������ڄ�������� ��܌��� ��܌����������Ώ�� ��������������Ώ������ Ҏ܎�������������ؙ�� Ҏ܎��������������ؙ�� Ҏ܎������ ������������ؙ�� ��������������ؙ�� ����� ӛ���� ��ȕ��� ��ȕ��� ������ؙ ��Ќ������������ ��Ќ�������� ��Ќ�������� ��Ќ�������� Ĝ����� ��̠Р����إ�������Ħ��������Ȩ���� ֤֤ؤ�� Ħ������ �������� ���Ȩݨ ���Ȩݨ ����������ƫ�Ӭج��Į����دۯ����������������° ͳڿ�������������������� Ѵ����ػ����ڿ������������ Ѵ����ػ����ڿ�������� Ѵ������ƺ�������� ̵��� ���������������������������� �������������������� ������������ ������������ �������� ����������� ���������� �������� �������� ������������ ������������ �������� �������� �������� �������� �������� ���������������� ���������������� ���������������� ���������������� �������� ������������������������ ������������ ������������ �������� �������� �������� ������������ �������� �������� �         ���� ������ ������ ��	�	� ���� ���� ���� ���� ���� �!�!�!�" �"�"�"�" �%�&�&�' �+�+�+�+ �+�+�+�+ �,�-�.�.�.�. �/�/�0�0 �
        �������� ������ ���������� �������� ������ ���� ���� ������ ������������ ������������ ���� ���� ���� ���� ���	�
�� �����	�
 �����	�
 �	�	�� ��	�� ���� ������ ������ �	�	�� �
����� �
�
�
�
�
�
 �
�
�� �������� ���� ���������� �������������� ���� ���� ���� �������� ������ ������ ���� ���� ���� ���� ���� ���� �$�%�%�& �'�'�'�( �)�)�)�*�*�+�+�+ �)�*�*�*�+�+ �)�)�*�* �+�,�,�,�,�, �+�,�,�,�,�, �/�/�/�/�0�0 �/�/�/�/�0�0 �0�0�0�0�1�1�1�2 �0�0�1�1�1�2 �0�0�1�1 �4�4�8�8 �4�5�=�= �5�8�8�9�9�:�D�D�J�N�S�S�U�Y�^�^�a�d�e�f�h�i�j�j�k�l�m�n�n�p �5�5�8�9 �5�6�9�9 �6�7�9�9 �6�6�9�9 �7�7�9�9�D�D�S�S �7�7�7�7�9�9�D�D�S�S �9�9�9�: �J�K�U�U�U�U �K�K�M�M �K�L�M�M �L�M�M�M �M�M�M�N �U�U�U�Y�^�^�a�d�e�f�h�i�j�j�k�l�m�n�n�p �U�U�a�a�a�a �U�U�a�a�a�a �U�V�a�a �V�V�a�a �V�V�X�X �V�V�X�X �W�X�k�k �X�Y�e�e �Y�Y�e�f �a�a�a�b �b�b�b�b �b�b�b�c �c�c�c�c �c�c�c�c �c�c�c�d �d�d�d�d �j�j�k�k�n�n�n�o �k�k�m�m �o�p�p�p �o�o�o�p�p�p�p�p �8�8�C�C�N�N �8�8�C�D �:�;�I�I �;�=�I�I�S�T �;�<�I�I �<�<�S�T �=�=�O�S�Z�[ �O�P�[�[ �P�P�Z�[ �P�P�Q�R�R�S �P�P�Q�Q�R�R �R�R�R�S �R�R�S�S �=�=�E�I�I�J�N�O�S�S�T�T�\�\ �=�=�G�G�I�I�J�J�\�\ �E�E�\�\ �E�E�\�\ �E�E�F�G�G�I�I�J�N�O�S�S�T�T �F�F�G�G�G�G�O�O �F�F�H�H�T�T �F�G�O�O�O�O �O�O�O�O �G�G�G�G�G�G�J�J�N�O�O�O �H�H�H�H �H�H�I�J�N�N�O�O �H�H�S�S �H�I�S�S �N�N�T�T �N�N�T�T �E�F�J�J �=�=�=�= �=�>�>�> �>�>�>�> �>�>�>�> �?�?�S�S �?�?�?�?�S�S �?�?�T�T�[�[ �?�?�^�a�j�k �?�?�^�_�j�k �_�_�`�a �_�_�`�` �?�@�T�T�Y�Z�f�f �@�@�U�U�\�\ �@�@�l�m �@�@�l�l�l�m �@�@�m�m �l�l�m�m �@�@�]�]�n�n �@�A�]�]�e�e�f�f�n�n �A�A�A�A �A�A�A�A �B�B�B�B �B�C�C�C�f�f�j�j �B�C�f�f �D�D�[�\ �O�O�Z�Z �T�U�[�[ �U�U�e�e �U�U�\�\�]�]�e�e �Y�Y�Y�Y �Y�Y�Y�Y�f�f �Z�Z�]�^ �Z�Z�]�] �\�]�]�] �]�]�d�e �f�g�g�h�i�j �q�q�{�{ �q�t�t�{�{�{ �q�r�r�r�t�t �r�r�r�r �r�r�s�s �s�s�s�s �s�t�z�{ �s�s�z�{ �t�t�z�z �t�t�u�u �u�u�u�u �u�u�u�u �u�u�v�v �v�v�v�v �v�v�v�v �v�v�v�w �w�w�w�w �w�w�w�w �w�w�w�x �x�x�x�x �x�x�x�x �x�x�x�x �y�y�y�y �y�z�{�{ �z�z�{�{ �{�{�� �|�|�� �|���Ӏ��� �|�}��Ӏ �}�}��� �}�}�}�~ �~����� ����Ӏ� ��Ԃ؂؂���� [    7   �          K   T   =   =   g   8     �Y<	�<4 t	=<4 t	=	K << f <P/< !  < < .<JJT��YO1 J! f J � J� , �J�X !@��~fY�����t�^��}JX�FX@g� y<Z�!x�� �"���v��~t !s �"���!}�3�X@/��2�  ���!q�;�X@/rv�J��!@�[Yos^��X!o �"���y�5rvWY�~���!@�[Yos^��X!q �"���}�XvF �Z�!~���f "(��X!� �"���x�6y$Y^�f��!� �"��	�!~�\Yu�Y
Xk�X!� �"����s�X��0/#�~\f}� *�!z�� y�"���!��XY$W[�f 0�!�x� "(�!��'�X@/#�6� !@���X@O� !@�Q���!@�[Yos^�� �Z�!8��~������~� !r ��!p�W^$Y��X@W�b\U[�~t "(��!�O���!@�[s���!@�[Yos^X� RP�4=f��gfuJ=u f=�$�=$�=��?? � � <5 � �1	�i	 h$ x�D �'�fN MX5 uX? H�s� ?  . f(     .M�	 �	�	=   <! �"     . J	K   "  . �( <.  <8 <;  * f .  . �<. F/     .  � < Y .( ..  <8 <;  * f .  .,�<�	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 �0 �- ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 �5 �2 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	��	=<f	�!  � <I' N3 - < ., !  f  K==<Y<, t> 2 < ., !  t	2XX*E�<, t> 2 < . X. /     .  J < K .( �.  <8 .;  * f .  .	�2�J+ a6 7� c� / T f\ 5 �8 �f �4 f�6 � �5 �7 � �5 �7 �6 �5 �6 �5 z�7 � �5 �: �8 �7 �5 �8 	�7 �< �; �9 �6 �7 	� ��@.<	-Y	Y<).f	/.�Z! Xm wJ	g�	z<f<-m. J�.20�	 �
J wX	 ��	 �G	 �K	 �K	 �K	 �K	 �K	 � �2 y	X 3 x. � � �2 � � X9�X�	 �/ J7X JJ	 ��	 �	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 �, �) ��	 �( �% ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	 ��	�0 M� �/ 6X / K.5X , O.. �/ �- � � � � � � � �, �. �- � � �0 �1  �0 �2 � �5 �1 �0 �2 � �/ �. �1 � �/ � �0 �1 �5 �. �/ �, �K �O �3 �1 �0 �/ �0 � �- � � �+��g	f�?�
  i�	=�	q.;�	Yv	K	K�	��	���	�<% m    ��	�g��(&���&)�	ef	��.3t�	g�-�<��"f	�#	�#X	<�	�=�%	�
  ��D � � �) z f f	� X	�"	1<�. �	�u�~<�����	-��~t ����>f�"*���"f��	#<% m ;Y��ffY0. � �	f	>�<f&U=�*8F��\X<	��$f < �D  <5&$.	q	�	��t	�J	��%	��K4 �=J �<	�#* S f f	= �	�"	h. �	�(�	[fZu��	f+ t �X�& x�u�(6�.t�.cf�~.Xf)�7����/&�( �v�f'<f��F+<X	�~4�x�hf�
� � � X 	�X�|f�1�%.=��1!< �!	u�!	�i	f	K$�|g	�*f	���| ��	g	� 	f�t	[���g#�t	�| 	���xX�4zJ( � �	��  K�"   I . �	M	Z   0  . J) J*    [0 I �Y"   ; . J	M	�  	#� tK�}  J X � fh��t7 �~X8   	{	Z|	�O �N�}  J X �	u�	� � �� �M �K�}   X �uY( �9 ' �8 �Y �K <�$� �K"I   � � � �K'Q �$ �4 x�1 ��$� �K <2 JA � �� <2 �D � �8 JG ��}  .$ �� �� <2 �G y� �7 JF ��}  .' �� �� <2 �E w�N �
<�}  .% �� �� <2 �F � � �K�}   X  �� �K�}   X# �� �K�}   X! �� �K�}   X" �� �� �K�|   X" �� �K�|   X! ��aLf5ff� �K#! �g��u �$ �&   Y J t�+ .-    X . �K�|   X% � �+ �| X�. �� ���|  J X ��) 	�= X��$�=&u'u%�K��w�. � �$ J&   Y ��"��Y   .+ �-     . J J .p�}  .& ����> < t# J J=@ < t% JuA < t& Ju? < t$ Jv�u. < teIJO<:<#<z�!	�U < t: J J# <=U < t: J$ t �YoiJJR<<<$<� "�^X�B<JJ$<=B<J%<�! �K�|   X! ��o� u  X"   /#! t�aLf5ffg ' X)    .! �Y �K�|   X" �� q�  X"    . �Y �K�|   X  ��o�#! t� ' X)    .  �Y �K�|   X  ��Y* �=  m�  .  J"    .* = �Y �K <4 JF l���|�� �8 �J � K�}	t �K	 �K	 �K	 �1 J � �3 �}. � �� �K <4 JF )L �BM �h ���}	t �K	5 � XK	 ��	 ��	 � � �� �K�|   X �� K�|	t �K	 ��	 ��	 �; J �# �� ��|	t �K	 ��	 ��	 ��	 ��	 �9 J �$ �� ���|	t ��	7 � X�	 ��	 ��	 ��	 ��	 � �  �� ��|	t ��	 ��	 ��	 ��	 ��	 ��	 ��	 �5 J � �� �K�}	t �K	1 � XK	 � � �� �K�|   X �� �K�|   X  �� �� <��|  .$ �; �M l� �� <K"$K�#5 �|�7 �4 �3 � �� .�"�$u#� �K�|   X �� �K�|   X �� �K�|   X �� �K�|   X �� �K�|   X �� �� u  X"    . e$ X&    .#! t� ' X)    .d$" tu   . �+ J-    .   X"    .e!*( tu     . �/ J1    .#! t� ' X)    .g! ��20 t J �   X"    .3 �|5 � ��&$ t� ' X)    .9 �| �3 v8 � �2 :5 � �3 ]5 � �: v � �  .  J"   /��{t) � J��" �33  	�	?(  ( . �	�; i< ,   , . J� JK u*:4.*rt�84 *r<*. J* f�>' X$ <KB�D*t<*.JJ*� ��/�<�=1$ t�� �~�t �~J	�� � M  f% �&     . JK�!  �C �!    fv�~��1�-Yu�K6<- �!/=;�-=*�XKf- ��6�7��~�	�*f	g� f.�7 K8   %X�J���~�[(ft~JM- _.    . JN?K%0?s�)! % ?;?. �$ J1 J? J`a�$�.$ ��(  $ ;$. JM�     J .I��~�� J �_��$�# � JH �6 fL,��%��~:�J�$��~��xJ	.,�1,<F ���~�J�1'!���)�*f��'$* *t> � t* �2"�%]�.lJ .5 �� ��k �s V  $ V .K J�"�K!  F J$�(' L �$�($(' K J$�(' N J$�(' O J$�(' N J$�(' M J �*K *. J;��~�I�	�*f	�f��-` BXh $   tY p<-XX	�	g� f.�4 J�"�K!%$<6 �)�J  )tJ . �_ Jg J  , J .6 J%K)7K(<)���<q.!Xu5!$6$i(' L �!�2J!�"2J!�X	�~	���.G LhG> , ��7 % � �A;%=6 , ;:6 0M �U 6  , 6 . J%K).7/(<)� t�%>(4 �<    X!2t!B2J!>2J!��%$ �%�>!�2t!���y !�.2J<��2��� [`t�g	g< t	Na J X.	rXY�." i<��.)�  	j.	�*f	�Y	�P�X� [�� <J��}��1*�.=��Kf��f&�&�,����P@6 J 6 .! �	���W �_ B   B <	KJ	��	K �2 J� �8 �� 7 J� : J� ; J� : J� 9 J �M�8J��}I�	�*f	�f��L B�T   	yJ	��	K<" ��6 <t6 . �K JS 6   6 <" JK#K<����
 8 ��<Z"<�^$�\'="  ':" 09 �A "   " < JK.#/<� t�f(  X XJ�L	h<J	�	�	u� t<k Jk<X	(�u�J<	�}	��	�J	�� t<m J�� ��*)t���x �� .����	�,2x�Ktu"0!�v	� <
 �	M� ��� <�		.
 �� J�`��G9<Y.*f ZX ���e<% J\<G,Y"�A?< J- �	�
 �X;��!�!K."�Ydt�x<�1-� .t�V*<��($f Jf!�N�,Y!j�!<f	=؂  �J!�".x��%� &tu�<JK�!��� <!KjX,Y��!C�� �,YJY!��% �j%	� �
 �
� .qX!��� <<AX%�j<< �tK	f�= �h�p
 	�$ �! �& �  �������x1��� �g�����	�	gJ	>Y�}����	q���	�}�x��})) �6	�tf�~�#��	�}J.Yg����*f<uw�K� �.!t<� <f$ � � �-P�.$ 7�( H  � /�Q K8 �& f�dD����6Xf) �K-�HL./<$��J<4 �� �$t;�V�� $�:� f�$K%�*i�5C�$t�%� c$ J�*�!) Jt�<G /( O.  � J	�f�f�!  f�g �Z$f��4f#Y�~�� 3~�gKM�*f<Kx3�<����$f�@�"'3#f Kg"X�=� = �)�"�1&�9X?��[��~8 �& f   �	�	��pf
 	cYZ	=	�.K/& y.   ��X<tX=f��g ���f# �. v	�fY	v$)t�	g)�	��)t	.�*f( �	�&�	��.	f& 	�L9Rt9.�}���Ngi�����4�4u$[&fK%fKJ<���f �~ 5 f �	���})��pJK�)��p�.f���1V�0 e�P��$<�?*t.*z��)fi	�!f* J1�2��fg2 t�fKC �~��*+>/f�><,��L3 f!=T!�'%!='!=+!�,!uA2f!�/t!����	�p"<f�����	�/&�	�� &.	���~ ��$f�@�$������ u"� �&�7�=��$f�[j��kJk�[t1,u<K-�.!./�X$�~�P<u@*t.*s��2�1���~��� @�$���� �g� �"� �&��9X?�$f�@�$���� �g� �"� �&��Xt�q.	�f�K$f��SX@��&<.,��&K��f� u"� �&�9�EX.X+&�f	�� �	g.	f� �<� �KfXj�g	 < t	 ��J �h�U�	 <u	 <�	 <�	 <�	 <�	 <�	 < �d-g��	wt1.un  �    u       < f��`.	
Jr. J   �J	)�=g  �    Y         <g<f�e=�%<�/<<�x.?��f	K	u6<	��Z�%ft	K	u6<	��h�f���f�	>	�	g"	�$	u"	�'	�	�	�	�	�	�	f��Y ��	'	"	gt-�	�g,.	t	�	�	�	��	�	�n�$ �!  & �  ����o"<f��������Y0<f<�E�N�f t	L, < �/4 W,    f		g�&?At2XYt<fY- f9 - <8? �- �fg	<�g]X� �g� ��� ���� ��=��f	�	u� �gsnt�!f	�	u � �" o. ��! � �u0 W    �	%	Y	u	Y�8g/ G ; < f(�t!Y<f��(�f& X� � V�0 X	�<�<�<�fY�	�)�	Y �Y$f/. J <H; Z.K<1 z�   fJt.	�J	>X/ J) <	��&�t7 J+ Y7 + < � ��= �+ ��!f/ JG ; <�>J# �,�m% /� ;��  � �  �f@ �/ g9     . �K ( 	<R  R � fg Jo R   R . J � �0	/� �=*���	��=	�- .	K& = �G &   J	ZL��		=�Y#	[J	! 	=.�����n#�K�<� 1u�	�mX	�?	��=	����X( 	�m� �J=	�� � ( �9 �J ���J.f �- .<# JY?(X�4r<4<! �4 ��3 <�2( �J ��  �mJ�@  �	�	�?�XE	 �=	�4	Lf� " /3 f=     . J	K%J=	� f=	Z	K�	g.���: lT �	� �@  �	�	�?tX) ?A �7 <��+ "-�!=$/� <A XP E <1 ,+  J X .X�*yXJ*u!< "T4%<F X[ J < ."/4%<F X[ J < .,�<Y	h���
 	& � 	& � 	& � 	& � 	& � 	& � 	& � 	& � 	%	=	u	�$ � ����rf�1�!!g< �h1���YY�����������f��1 �r< �    <   �          �   �   z   z   g   �   @ 0}  g	 "     	Y.< J& * <1I/;h! ��K�g	  X.! �  	�f � �t& yX5'��	�	K
 s4!./��	h�����f�/I	r. J . J� qJJ@���Y<f&J�K .�g+h�	 t# f  	u u�" J" p X9�i]^ J�r;<X��	sf�<nf	
�D7k� ' �/ # <   J <+ J/=  	-.=  )7 ���x'��	!<P	��X	/	�	�u>!f�(�11<-h8) - 1I1. J1 X['<�<K��fN�-�<h�"/ ��Ju�!{Y�: $ : < � : t�CG : I$ : J* � �w< $ < < �K?C < I$ < J+ �< � �	J<P2�Y�!�tg�#%1�
�	[<S	�	�	�#	�  �1 	>!	�	�K	��.	�	�#	� �0 	?!	!	�<.�1J��y<z�2. i .�A<  ,;�!	 �# �  	�&tf �7 t> �Js/5��. �K �� f. tv� ��!�"/{L��f��	s�;  S �	�	fgx<.	l�<	f�'�!	f JKf	KL\Xgf J <  J J JK  = |=gf J <  J J JK  = <!�	f�@)��"L	 ���	t<	� �	�2	zd<0 J�= b  �Y,�/J.K+�)� cf J J !v��f�j���g�?Jf< � � � ff�f�<fgf�h���u� J�� t�� t��!uu z� � ���!K� t  f J �= ;KL!	 �s�- � <9 �   + . J
Z%Zu }+ .g J t	�&	Y &-.0<�� t9 t ��)� ��Y�L�' J�K �/ t J, <	u��	| Xu%� � yf/f% t�
f	s�f+ J�%� �h. �	m�8��M<t�t	g��<B��� � f��|��|�	 �.��|��|�	 �.x�M'����J�J$�&	u	I[����
 �E . � J	�w:�	�) pX J J <	�	�	���@X�	@2E� � �	�	���#��('*"� � f���0 O� .�+ ��� .5��� J�;OY�L�{��{�.��{� J fH�{�." �6 f, fi< � <( J" <: f0 <	gYF );XN�t	s[$  f	F( @G f8 .	gfX	[f .��*iS t4 <�.Vft��	if2 J f7 JO �C f	g	gjf1 � X6 �N �B f9 c� �0 s
�0<��E<tf'���LyyxfX	p�u	]<f	��t, XY-�-�	p	g. J: 
 �V    <   �          �   �   �   �   �   �   1 D�  �!   . �$ J% )  *  <  . f .K.Y;<.Y-5�~J�f�:<f��
 	� ; 	 I  t� =�JtJ		��f �  �.� .f �. X       <K<	� �� .+�X�Ep<<D	�	mY.�	 Xs�&K	�<	m�� ���	� 	�	Y� �	�~��	=�0 
Z+ � <�&J/��h&=J	�d<g&g	�<e z�#  d� .&
f=	\<f�Ue�k&Y	xf<1g�J1 k&Y	u	��	�teւb&g	�ft		�X<g&g	�	��� I�<v��� �_J  <�J ���IJ	� 	��. Ys�~KX� I= I �� D	� �	Z�
 � � �. � / J f( J) -  .     . � . J#   < < � JM�		��= 5I �� ��	�$ �   .J��~&
�/	�:< �KY��~�&
JK	�H< �  �� �� �	T	��<� f- 2� J8 $<�< .K� &
�K	\d< � r��	� 	Y	uJ>��	�~J	=t	=�� �&
�.K	N:<	� 	�*�� �.�J��* � !�&
f/	N<f� �J�J. � � X*v�"� J	�J	K�	=t�  t*v�X	� 	YX� Kg' ;  &K<' ;   J � J& � � �X J . �$ J% )  *    / - J J, �  & < <�JJ � K���}  � �       <g<�' 3 f�~u&g	x</ �'  �~�<3 ��~�		=�	� 	YXt X*v�X	J	K�� 	J	Y( ��&g	x<	� uX�&
f/	Nf� "�.f	J	Y 	��	=�"� .Y.	�X	=t� "/3��fw�	J0+��f	K	��tyf	Jt3�}J�	Kh."�	Kh<"�	K	g'�>;>�	K	gvC0Y�	K	h�~<  �       <g<��.�H JH ��K �K ���~   f � . �$ �% )  *    = - JK �	� J	X�! 0�/<K ��tH W <J^)�|<  t f       <g<� � �� �3  �~� �$ J% )  *    = - � J $ J% )  *    = - JK � �~J $ J% )  *    = - JK � J!  J J � ,<�~� � �!  � u!  � �~� �$ J% )  *    = - JK � J!  J J �hX�Y�!
�#�|J  �    u       <g<X � $ �% )  *    = - JK �	� �	�.	�#i*" .�J�.�|�  �    Y t �       < ��../�J�!J0 +�%Xu�<2��X� �~� �$ J% )  *    = - JK � �~� �$ J% )  *    / ; JK �	� �	�.	�#1* bf*  � % "$eQ��~<  =t ; f$ J% )  *  <  . f .K) ��~<�<.�� z�%   �~�$ J% )  *    / - JK ��	 ��	 ��	 ��	 �	 	KO � .W Xw �	�R! � �[ X| X	/�R Ǟ.	 �	KO J .W Xw X	�R! � �[ X| X	/�R Ǟ.� p�"  f �"  !  f �!  f"z�fR�A<) X0�}���	K	hfY7 �=�~
 	g ; 	 I  < J�/v��	K	hfY5��=�~
 	g ; 	 I  < J�&hK	Kh(0K J ��	hB�.YL!!(X�\c�#Xd�& t f�<f�=YK
�*<J�x��_& d�	�K��J ).$���<2J �# �BJYL.�m��o��Xr�=   < f      .KK.91" I0&tf=.� J .�A v�' ( =<( s" .�CJ!L.of�wt�5tX�Xyf^�� �: �- < �  f �x���	u)�z.   . �$ J% )  *  <  . f . J2 �  {<	Y=�x�  �       <g<	�":f	�v�z�< �)K<)�K	 �z� fR��� J: X- < P  ff	u)�z.   . �$ J% )  *  <  . f . J2 �   t	.�z�< �)KJ)�f�z.M�fK J9 X, <Lf	Y&*�vK"/ J9 X, <N �	�
�	b<;^K J9 X, <KH �0#4�w
 	� ; 	 I  <�JHJ�fZD��wf  f       <g<�=���/< vJ XBX��z
   f�	K�   . �$ J% )  *  <  . f . J0 �    t�/�y�< �  J�  >.�y<N���
   f �w���	�&�y.   . �$ J% )  *  <  . f . J0 �  {J	Y8�w�  �       <g<	�5f	�;	�v�yt< �&KJ&tu
 �yf f/���*>K�u9B�u;h���E$�uhG��uh4�z���~f�<J�<��� �f$X� ��}	�	���	���{�  � �       <g<	��~	�	�	��}	�v	�<	��}f
   f�f	��   .  $ J% )  *  <  . � . J0 �    � 	  f��� �	��   .  $ J% )  *  <  . � . J2 �    �	��	�}��t�<���f	��~�	vXy	�	��}X�< �  �	�  � t��|<< � ���	/g*f #J=�	�~�~t   J �$ �% )  *    / - JK ���~	�	��\�X�	� �|�   J �$ �% )  *    / - JK ���}	�	��"��}f�� �|�  t � �$ �% )  *    / -K+ � ��}�		�	vX � .$ J% )  *    / - JK � �~�  $ J% )  *    / - JK � �~�  $ J% )  *    / - JK � �~� �$ �% )  *    / - JK ���~	�	���~	�zf� �{�<	��}  � $ J% )  *    / - � J  �$ J% )  *  J J / - � J .  �  �$ �% )  *    / -K ���~	�	��� .��f �}J �$ J% )  *    / - JK � �|�  $ J% )  *    / - JK � �|� �$ J% )  *    / - JK � �|� �$ �% )  *    / -K ���}	�	��#uW J��	�}	�	� ��^�	�} 	�	�1<<�f��| ���~	�	�����}	�	��Y�}f.����. �|�  t �$ J% )  *    / - � J��}M�<z��1< �zX t       <g�<�}	�	���}	�i�<��}	�zf�< �z� < � �  �  �$ �% )  *    / -K/ ���}	�	���}	��t�}<fX	vXy	vX �  t � <$ J% )  *    / - � J��}J�. ���}�	vX �  � � J J$ J% )  *    / - � J f*� �}�  < � �$ �% )  *    / -K* ���}	�	����}	Z�< �z�     Y    X��z      Y �       <g<��}	�	����}	X��}�	X��}X	X��}�	���	vX�/ ���}	�	��'ut�}f� �  t ���}�	tufX��~	�	�����}	�	��Y�}����}�.� �|� �$ J% )  *    / - JK. ��$uK�}� �|f  � t �$ �% )  *    / -K/ ���}	�	���}	KX�	�}��	���}�	���}f����}	���~f� � �	� � �} ��	vX� ���~	�	���~	�v� �}�J�~�f	��}  ' ��� �}� � �  �$ �% )  *    / -K ���}	�	���}	t � X	�  t	u�}�	�	�&y� �|�  f J J$ J% )  *    / -K& � �|J  . f$ J% )  *    / - JK# �	��|	�	�	x� �  t � �$ �% )  *    / -K' ���}	�	���|	� �J �$ J% )  *    / - JK' � �~� $ J% )  *    / - � J  t��}	�	��#uY' J . ����}	vX	t�	vX�y	���~.	vX	tz�	vX�. ���~	K	���~	�v� �}�<�~�f	��}  �� 	���~�	vX�<W�X&��|   t � . t$ �)    t! � JK �	�� �z . f       <g<��~	�	��%Y�~���#ff�_�"�{  �       <g<� f�&�	�~X�J	vXy	t��}.	 �t� t��|  � t  �$ J)    t! � JK% � �|� t$ f% )  *    / ; J fK � �|� t$ f% )  *    / ; J fK � �|� $ J% )  *     . J .K � �|� $ J% )  *     . J .K � �|� $ J% )  *     . J .K � �|J $ J% )  *     . J .K �	�� �| � . �$ J% )  *    / - JK+ ��~�� � �$ J% )  *    / - JK+ ��~��	t��|<�D � �~� �� 	vXy	vX�u)�.Y�&Y+ u+ -V ��+ yt
.u; �1 <. ��u"-���"�~.< mX2 </ ���	�	�	�	� �|/$ J% )  *     . J .K �	� J t		X�9�~���XX�=0/<K<��B<W-X �|  < f$ J% )  *    / - JK/ ��u� �{X t � ��	vX �� �$ �% )  *     . .K �	�k � f��~uv& K#&�~��j/$�/ -Z Y=���#rJg u-��~f	K� �  < .$ J% )  *    / - JK3 ���� �} J$ J% )  *     . .K �	Kw	f � f��|f	��}  X	��	t< f	K J J	���|
  �	�(�.(�  �� J   �  t � � t�J � 2 �   .	���{J � 2 e   . �. ( �! f	�7�u��|��	/	��{   J . X$ J% )  *    / - JK � �{� �$ J% )  *    / - � J   $ J% )  *    / - JK � �{� �$ J% )  *    / - JK2 � �{� �$ J% )  *    / - JKF � �{� �$ �% )  *    / - JK ���|	�	=��!u XK�|���,���{< �}�|	�	�  � �$ J% )  *    / - JK � �{� �$ J% )  *    / - JK0 � �{� �$ J% )  *    / - JKC � �{� �$ J% )  *    / - JKV � �{� �$ J% )  *    / - JK � �{� �$ J% )  *    / - JK1 � �{� �$ J% )  *    / - JKF � �{� �$ J% )  *    / - JK � �{� �$ J% )  *    / - JK3 � �{� �$ J% )  *    / - JK � �{� �$ J% )  *    / - JK0 � �{� �$ J% )  *    / - JKD � �{� �$ J% )  *    / - JKX � �{� �$ J% )  *    / - JK � �{X$ J% )  *    / - J J ��.Y$�.Y8 �. <+ ��u)uW( �! . �( � �	�|�	�X	t�<	hXU � J=( J�6
Xg�|f��f��{����0 i.�{t   <   J$ J% )  *    / -K# �	K�|	�	=�	�	!�|	� �{ �*�*<Y���|	���*�*< �{X  f   J$ J% )  *    / -K* �	O �{  . < �$ �% )  *    / -K' ���|	�	�	x�	���0 ��{<   < J �$ �% )  *    / -K# �	��{	�	��	�Xy	hX	t�J	v<��#u���yu��~ 	 / t    g �u������z<J���zJ/ �	�	�/��z	��/ ��?� ����/�=g�v��v��u ELEM_BUTTON ELEM_FIGCAPTION visibility attrs_len close fs_rename PARSE_DOCTYPE in_script size_str cursor_move_right border_bottom strncmp tab_title parse_flex_wrap ELEM_FOOTER cursor_move_end nav_home tag_name rel_len mem_used block_y_start version dom_append_child ELEM_HTML kernel_api_t input_cb_t cache_find element_type_t layout_computed history_entry_t first_child text_run_count ELEM_LI content_margin cursor_backspace ELEM_PRE parse_position handle_end_tag fetch_url ELEM_TH link_x word_len attr_ptr style_str border_top ping font_size text_w class_name exec extract_origin margin_top search_mode parse_overflow ELEM_ASIDE is_auto active get_fs_generation oldest tab_width text_run_t send scheme_len ELEM_TITLE uint32_t fg_color ELEM_SCRIPT page_title fs_read scroll_offset vals PARSE_DATA page_content memmove current_padding_top malloc cursor_x str_casecmp nav_forward cache_add box_shadow_x box_shadow_y scroll_h result has_border fs_exists long long unsigned int browser_tab_t strncpy content_width lib_name border_width margin_left parse_align_items parse_flex_direction has_content parse_size ELEM_HEADER box_idx ELEM_FIGURE parse_align_self current_tab encoded write_content extracted box_shadow_color ELEM_OL block_stack draw_text_clipped execute_script_content dom_node on_paint css_style_t block_x_start toolbar_y tag_len total_height z_index next_sibling history_pos open_url_new_tab set_window_menu copy_len url_cursor_blink q_param block_x free current_url recvfrom link_url font_weight text_start dom_node_t draw_border flex_shrink line_height mem_total DOM_TEXT ELEM_TEXTAREA type_attr ELEM_SPAN win_handle_t base_url menu_cb_t fs_delete nav_back font_style page_offset tabs PARSE_TAG_CLOSE border_radius dns_resolve dom_create_node border_right ELEM_LINK parse_border_style exit ELEM_TABLE switch_tab http_get flex_grow url_encode parse_html action_id ELEM_BR name_start dom_nodes ELEM_OPTION target_blank page_cache_t entry max_width extract_google_redirect host_end str_cat long long int ELEM_A ELEM_B ELEM_MAIN cdl_main ELEM_STYLE valid ELEM_I page_cache ELEM_STRONG slot is_loading href ELEM_P html_len text_len ELEM_DIV ELEM_U PARSE_SCRIPT ELEM_BODY link_y write_len parse_color fs_list target value_start itoa scroll_pos exec_with_args content_w history border_color current_element dom_node_count max_chars max_len cursor_move_left cdl_exports_t text_runs handle_start_tag default_style paint_cb_t GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection border_left content_height tab_x path_len ELEM_SELECT centering_offset color_str ELEM_SECTION text_decoration get_element_style ELEM_TD box_run_t draw_rect sprintf parse_justify_content parse_state_t ELEM_TR origin_len DOM_DOCUMENT symbols elem_width item_count unsigned char PARSE_ATTR_NAME print script_buffer_len ELEM_TBODY ELEM_HEAD parent short int get_kbd_state connect history_count final_url display draw_rounded_rect get_launch_args style_attr loading_dots quote PARSE_TAG_NAME attrs ELEM_UL max_text_width ELEM_EM fs_create title_len PARSE_TAG_OPEN tab_bg draw_text list_type block_h value_len val_len link_region_t cached block_w min_width block_y on_input create_window socket has_background draw_rect_rounded url_cursor_pos content_y res_len text_align fs_write process_events DOM_COMMENT padding_right on_mouse box_shadow_blur ELEM_DETAILS cdl_symbol_t prop_len resolved_url sendto tab_bar_height is_url ELEM_LABEL elem_type box_run_count is_link text_buffer bind list_counter parse_state prop symbol_count ELEM_META navigate bg_color is_closing ELEM_SUMMARY script_buffer skip_depth ELEM_H1 ELEM_H2 ELEM_H3 ELEM_H4 ELEM_H5 ELEM_H6 ELEM_UNKNOWN func_ptr word_start text_node DOM_ELEMENT ELEM_BLOCKQUOTE ELEM_HR ELEM_IMG layout_dom draw_x draw_y margin_right draw_image_scaled relative_url current_padding_left mouse_cb_t net_get_interface_info label resolved PARSE_COMMENT link_region_count realloc timestamp alt_len ELEM_ARTICLE content_len recv content_h execute_document_write padding_bottom cache_restore short unsigned int dom_node_type_t block_stack_top cursor_move_home memcpy flex_basis last_child ELEM_FORM ELEM_INPUT display_text status last_slash ELEM_THEAD add_box_run ELEM_CODE PARSE_ATTR_VALUE margin_bottom resolve_url aligned_x link_regions ELEM_NAV box_runs get_ticks cache_count handle_text tag_name_len tab_count tab_index cursor_insert_char text_content menu_def_t parse_inline_style max_x scheme_end strcmp get_element_type key_content_end hlen cm_bind_action clist_path parse_plist_xml file_buf my_memcmp my_strchr cm_dialog_select_dir file_picker_cb_t perm visible_items start_dir cm_dialog_submit show dates my_strstr parse_menus_from_string cm_dialog_input selected_index config_count current_dir cm_dialog_save entry_count val_tag name_ptr full_path initialized real_idx nlen default_name menu_end key_tag i_idx cm_dialog_handle_mouse dirname max_read file_picker_t cm_init temp_menu_count cm_dialog_open needle temp_menus action_bind_t execute_action_by_id entries strncpy_safe cm_dialog_click filename id_p req_h haystack menu_idx cm_picker menu_tag req_w cm_dialog_up_dir cm_get_config list_h cm_picker_refresh list_y is_dir item_h buff klen config_pair_t key_content_start icon lbl_p action_count cm_dialog_render cm_dialog_init cm_apply_menus func val_content_start vlen cm_load_app_config item_tag cm_draw_image_clipped win_handle win_h flen win_w win_y filter filter_ext val_content_end item_ptr key_name raw_entry_t internal_menu_callback filename_input app_bundle_path win_x cm_draw_image item_idx actions safe_div2 body local_count keywords is_alnum js_set_global dom_window js_console_error js_console_log js_to_number TOK_PUNCTUATOR TOK_ERROR condition values js_window_setInterval js_get_global this_value js_strlen functions next js_value js_get_error TOK_STRING cond js_new_string function_count is_keyword JS_TYPE_OBJECT number_value init_lexer js_strcpy js_new_undefined next_char js_array_length js_strcat skip_whitespace TOK_NUMBER js_array_get js_value_data_t js_property_t function_id js_array_t js_new_array parse_expression heap_used column locals js_new_number js_object_set parse_function_call elem js_window_alert js_register_dom_api operand param_count parse_primary operators data js_type_t js_array JS_TYPE_STRING property_count js_value_t error_msg call_stack js_new_object js_clear_error TOK_IDENTIFIER parser return_address TOK_EOF JS_TYPE_NUMBER js_object_get js_object_t has_peek source numbuf js_function_t js_value_unref console next_token elements JS_TYPE_UNDEFINED token_type_t js_console_warn js_to_boolean cond_true js_call_frame_t engine current js_variable_t js_document_querySelectorAll is_alpha static_objects is_digit js_eval lexer_t dom_document find_variable scope_level js_memset is_native js_new_null false_val parse_statement eval_binary_op str_eq prototype js_init JS_TYPE_BOOLEAN js_to_string native_fn token_t JS_TYPE_NULL properties js_engine_t heap js_document_querySelector advance_token params js_window_setTimeout obj_idx JS_TYPE_NATIVE_FUNCTION static_arrays js_document_getElementById line ref_count true_val has_error global_count find_function TOK_OPERATOR condition_start peek_char call_stack_top current_token uint8_t print_callback js_object JS_TYPE_FUNCTION TOK_KEYWORD js_register_native parser_t js_new_boolean argc arr_idx value_count alloc_value js_array_push globals JS_TYPE_ARRAY max_iterations js_value_ref /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/apps/browser_cdl.c usr/apps usr/apps/../../sys cdl_defs.h usr/lib/camel_framework.c usr/lib usr/lib/../../sys camel_framework.h usr/libs/js_engine.c usr/libs usr/libs/../../include types.h js_engine.h    ���� |�  <           c   A�A�A�B
�A�A�AI
�A�A�A  <       d   �  A�A�A�A�CP�
A�A�A�A�D T       d  _  A�A�A�A�C$
A�A�A�A�De
A�A�A�A�C   \       �  +  A�A�A�A�C0�
A�A�A�A�CF<G@K0Y
A�A�A�A�C $       �  p   A�|
�CR
�B[�        `     0       p    A�A�]
�A�D�
�A�A   <       x  �  A�A�b
�A�C�
�A�AF
�A�A   ,       4!  H  A�BI���:
�A�A�A�C �       |,  �  A�A�A�A�C0�4E8B<E@w0E4A8D<A@Z0m4G8D<G@J0C
A�A�A�A�AR4A8D<H@R0C
A�A�A�A�A   P       T.  �  A�A�A�A�F��
A�A�A�A�B��G�H�L�   x      C    A�A�A�A�F� J�(o�(A�(A�(P�(��(H�(b�(O�(A�(G�(U�(��(E�(B�(A�(|�(Q�(A�(D�(A�({�(
A�A�A�A�A�(E�(B�(E�(i�(B�(A�(I�(w�(��(A�(A�(A�(P�(H�(E�(A�(D�(C�(j�(B�(A�(P�(L�(F�(B�(A�(P�(P�(��(A�(A�(A�(P�(P
�(E�(A�(TA
�(B�(A�(TA�(B�(A�(P�(]�(g�(E�(A�(P�(P�(b
�(B�(A�(TX        N  �   A�A�A�K
�A�A�DP
�A�A�BU
�A�A�AM
�A�A�Ad      �N  D  A�A�A�A�F���E�B�E�k�B�A�I�B�
A�A�A�A�Dp�A�A�A�P�j�B�A�D�L�U�E�A�D�P�R�E�A�D�P�E�A�A�A�S�K�B�A�P�P�y
A�A�A�A�AA
�B�A�Q\
A�A�A�A�AA
�B�A�Ti
A�A�A�A�AA�B�A�P�]�r�E�A�P�P�X        U  "  A�A�A�A�F� J�$�
A�A�A�A�D\
A�A�A�A�D `      DX  �  A�A�A�A�F�\�G�G�m�T�G�A�F�_�G�K�J�E�B�G�s�E�B�G�F�E�A�G�O���D�d�N�D�f���D�G�J�H���A�U�i�D�A�E�J�A�G�M�����G�H�H�A�D�L�}�y�G�P�J�A�E�T�k�A�G�\�J�A�G�Z�F�O
A�A�A�A�A��G�D�J�h�E�P�L���D�I�L�L�G�G�}�A�G�A�J�A�G�\�J�A�A�Z�L�B�G�X�i�h�G�E�R�Y�G�V�g�A�D�B�R�f�G�V�g�A�D�B�J�b�G�G�A�b�A�M�D�F�         j  �  A�A�A�A�F�\
A�A�A�A�BC�G�A�L�G�A�A�L�K�A�E�L�C�A�]�F
A�A�A�A�DC�G�A�L�G�G�A�L�K�G�A�L�K�G�A�L�K�G�A�L�K�G�A�L�K�G�A�L�v�G�E�L�Y�G�A�L�  0       m  O   A�A�A_NG TAA�A�0       hm  V   A�A�AfNG TAA�A�,       �m  5   A�A�CXG NA�A�         �m  �   \�F F   t       �n  s  A�A�A�A�C0f8A<J@J<A8H<G@t0L
A�A�A�A�BY8A<E@L0U<A@H0F8G<A@0 �       p  �  A�A�A�A�C<V@O0c
A�A�A�A�AC<A@U0z
A�A�A�A�E{<A@H0c<A@_0\<A@W0@<A@Q0   0       �r  8   A�A�AWGF NA�A�   |      �r  W  A�A�A�A�F�u
A�A�A�A�AA�J�J�t
A�A�A�A�C��A�L���A�A�H�S�W�E�A�E�d�Y�A�S�C�A�S�T�A�S�D�U�J�D�C�P�T�E�A�A�X�h�A�K�V�X
�E�A�E�R]�E�J�E�M���A�L�@�E�A�H�S�m�A�A�E�]�D�Q�H�A�D�C�P�a
�E�D�E       Lz  �  A�A�A�A�C(\,F0t w(G,G0R g$E(B,A0R I(F,F0F4E8E<G@N(G,G0T,A(A,D0J,A(G,D0J,A(G,D0J,A(G,G0J,A(G,G0T,A(G,G0J,A(G,G0J,A(G,G0J,A(G,G0T,A(G,G0J,A(G,G0J,A(G,G0Q4B8A<A@HA�A�A�A�C ����       ��            ��            ��            ��            ��        ���� |�  ,     0}  5   A�A�k
�A�BC�A�   l     h}  �   A�A�A�A�C0^<D@O<D@O0a4A8D<A@H0K
A�A�A�A�CGA�A�A�A�        ~     D      ~  �   A�ClG EEBF @A�B�W
A�DCA�0     �~  N   A�A�AZJM VAA�A�X        |   A�A�A�A�C0|8D<A@L0W
A�A�A�A�ECA�A�A�A�T     �  �   A�Cl
A�CCW HC
A�BCG HC
A�BCG HCA�,     (�  8   A�A�k
�A�BF�A�   �     `�  �  A�A�A�A�CTaXB\K`NP}XD\A`NPKXD\A`JPgXK\A`LPAXD\A`NPiXG\A`JPGXK\A`JP�
A�A�A�A�A(     ��  �  A�BF�����A�A�A�X     ��  v   A�A�A�A�C0w8D<G@L0O
A�A�A�A�DEA�A�A�A��     0�  �  A�A�A�A�F�Y�e�A�A�E�Z�N�G�C�K�L�A�G�A�G�C�W�I�E�B�A�L�E�A�A�L�K�A�e�K
A�A�A�A�BC�G�m�H
A�A�A�A�AC�M�E�,     Ć  D   A�ClAGA FCA�       �  :   A�t
�CA�     D�  :   A�t
�CA��     ��  3  A�A�A�A�CLRPQ@_LEPH@IDEHBLAPLDBHALDPN@@HDLAPF@]HDLKPF@~HALTP[@bLAPo@C
A�A�A�A�DCLAP\@MHALJPL@  4     ��  V   A�A�CX EKBG ]A�A� d     �  �   A�A�A�A�C z(A,D0N G(A,D0N G(A,G0]A�A�A�A�B ����  D     Ċ  \   A�A�ASDDD U[
A�A�DAA�A�   X      �  �   A�A�A�A�C(R,J0L G,A0O m
A�A�A�A�AO(A,D0L  T     ȋ  {   A�A�A�NJ ONGC LLD GADC JA�A�A�   �     D�  �  A�A�A�A�F�j�D�E�]�R�G�E�L�G�E�C�L�J�G�O�P�A�G�A�A�C�K�G�A�E�L
A�A�A�A�D^
�A�I�A�P�C�DZ�H�J�M�G�A�L�       �  �  A�A�A�A�C@`HBLEPETEXE\I`FHBLEPETEXE\E`LLEPBTEXA\A`LLEPBTEXG\A`LLEPETBXA\A`LLEPETBXA\G`SHBLEPBTBXD\A`S@EDGHALHPNTDXA\H`LLEPETDXA\K`S@ZLBPATIXA\A`LLEPBTEXA\A`LLEPBTEXG\A`S@lHBLBPATHXA\B`H@EDQHDLHPW@eLEPBTEXD\H`L@JDGHALHPbTEXA\E`LLEPBTEXE\A`L@EDGHALHPL@GHBLEPBTBXA\O`V@EDGHALGPJLAHBLEPBTBXE\G`U@NDAHALJPE@H
A�A�A�A�CaA�A�A�A�     ��  %   T     ��  �  A�A�A�A�C0�
A�A�A�A�Dy4A8N<G@F0�<H@H0(     ��  �   A�Cs
A�DOM I      ��          ��          ��          ��          ��        ���� |�      �  D�  <   A�i
�BK
�A ,   �  ��  �   A�A�i
�A�Dr�A�  l   �  $�  f  A�A�A�A�F��
A�A�A�A�AK
A�A�A�A�A�
A�A�A�A�A  4   �  ��  @   A�A�F�U
A�A�A]A�A� @   �  ̝  [   A�A�A�F�l
A�A�A�D[A�A�A�   �  (�        �  <�        �  P�  "      �  t�        �  ��  4   A�r�   h  �  Ğ  )  A�A�A�A�F���K�D�J�F
A�A�A�A�B_�A�D�J�F
A�A�A�A�D��D�D�J�F
A�A�A�A�CK
�OC
�P��T�D�J���B�D�J��
�A�UO
�Oy
�JH�B�D�J�F
�A�O��A�A�D�J�o�A�A�D�J�T�D�J�F
�A�PA
�A�PA
�A�PA
�A�PS�A�   �  �  a   A�_�     �  T�  ^   A�\�     �  ��        �  Ħ  #   �   �  �  l  A�A�A�A�CPhXG\D`HPC
A�A�A�A�CCXG\D`HPC
A�A�A�A�CCXG\D`HPC
A�A�A�A�CPXA\D`HPC
A�A�A�A�DYXE\D`HPC
A�A�A�A�CC\A`HPE
A�A�A�A�C�   �  T�  �   A�A�A�A�C g(B,D0H C
A�A�A�A�AC(K,D0H C
A�A�A�A�CC,A0H E
A�A�A�A�CI(A,D0H C
A�A�A�A�C   �   �  P�  �   A�A�AiBD HA
A�A�CKBD HA
A�A�DCLD HA
A�A�BCA HC
A�A�CC   P   �  �  �   A�A�A�A�C�
A�A�A�A�C\
A�A�A�A�A\   �  �  �   A�A�A�A�C0f<D@L0C
A�A�A�A�DY
A�A�A�A�A      �  ��  0   (   �  ̫  Q   A�CvD HC
A�B    �   �        �  @�     ,   �  \�  �   A�A�A�|
�A�A�A H   �  �  k   A�A�A�A�I
�A�A�A�DK
�A�A�A�A P   �  T�  �   A�A�A�A�A�
A�A�A�A�BZ
A�A�A�A�A   �  H�  
      �  T�         �  l�     A�CM HA�  $   �  ��  !   A�COD HA�   $   �  ��  !   A�COD HA�       �  Ю     A�CM HA�      �  �     A�CM HA�      �  �     A�CM HA�      �  $�     A�CM HA�  �  �  @�  �  A�A�A�A�F�}�F�P�J
A�A�A�A�AL�A�P��
A�A�A�A�AV�A�H�p�B�F�P�J
A�A�A�A�A�
A�A�A�A�F�
�A�D^�F�F�P�J
A�A�A�A�A^�D�F�P�J
A�A�A�A�Ar�F�P�k�F�X���D�D�F�R�s
�B�Ef�F�P�d�A�D�F�L��
�A�E�H�A�P�R�F�P�e�A�H�A�P��F�P�a
A�A�A�A�Ef�A�H�A�P�F�A�H�A�P�F�A�H�A�P�F�A�H�A�P�
�A�B�ED
�A�A�F��A�G�A�P�V�F�P���A�G�A�P�Q�A�K�A�L�h�A�G�A�N�F�A�B�A�P�b�A�B�A�P�p�A�H�A�I�H   �  ��  T  A�A�A�A�F�z�A�Z�b
A�A�A�A�CH   �  �  �  A�A�A�A�F�L
A�A�A�A�Ba�F�L�H   �  ��    A�A�A�A�F�	��	A�	J�	rA�A�A�A�   $   �  ��     A�CMB HA�   $   �  �     A�CMB HA�   L   �  <�  c   A�A�CP HAGA PAGA PAGA HA�A�    �  ��        �  ��        �  ��        �  ��                                 ��       c        d   �    -    �  �     ;   `�  �     H   d  _    T   `I      b   �I  4    k   �  +    ~   �1      �   �  p     �   `       �   p      �   x  �    �   d�       �   � H	    �   �      �   l�      �   p�      �   �}        �}  �     |,  �    #  @�      -  `�      8  �5      G  �5  �   Q  d�      a  D�      s  `�       �  T.  �    �  C      �   N  �     �  �N  D    �   U  "    �  h�        �5      
  @% `      ��      '  (%      3  x�      A  `�       M  �� @    U  �� �g    b  j  �    w  t�      �  @�      �  �         �  �U         �  �l         �  Ll         �  \p         �           �  �         �  <         �            �  �         �  �         �            �  �         �           �  4         �  �         �  �	         �  �          �            �  �         �  h         �             �           �           �           �           �           d           t         $  h         )   	         .  �         3  
         8  P         =           B  �
         G  d         L  <         Q  0         V  �         [  �V         b  XV         i  �U         p  �U         w  �V         ~  8V         �  �U         �  m         �  pp         �  �p         �  �p         �  �p         �  Xq         �  pq         �  �q         �  �q         �  �q         �  �q         �  (r         �           ��~   `N      �  @J         DJ        `J                 ��'  D�  <     .  ��  �     :  $�  f    E   �  X     N  ��  �     X  ��  @     f  ̝  [     t  Ğ  )    �  ��      �  �o     �  �o      �  �N  !    �  @�  �    �  ��  T    �  �  �    �  �         �  T�         �  t�            ��           Ч           4�                      ��  ��        (  ��        >  ��      	 G  ��        ]  ��        s  ��        �  ��        �  ��        �  ��  !     �  ��  �    �   �       �  ��  �     �  <�         �         �  �    /  �G      <  ��  %     S  �~  N     b  �m  5     k  ��  4     y  T�       �  ̫  Q     �  P�  "     �  l�       �  (�  8     �  DX  �    �  �>      �   ~       �  P�  �     �  ��  3      �  :       @�        D�  �    ,  Ċ  \     ;  T�  �     H  hm  V     T   ~  �     \  H�  
     i  `�  �    �  ��       �  �r  W    �  ��       �  �  �     �  ��       �   �  �     �  p  �    �  Ħ  #     �  D�  :        (�         �  �        �  �     0  ��  v     >  �  a     L  T�  ^     Y  ��  �    i   H @    q  ��       }  $�       �  \�  �     �  �n  s    �  t�       �  h}  �     �     |     
  �m  �     �  0�  �    �  �1      �  m  O     �  4!  H    	  �       �  �>  	    !	  ��  ��    .	  Ю       I	  ��  0     W	  Lz  �    `	  <�  c     t	  �  k     �	  �  l    �	  ��      �	  ��  !     �	  �       �	  T�  �     �	  ��  V     �	  Ć  D     �	  ȋ  {     �	  0}  5     	
  @�       
  �r  8     "
  �  �     9
  �  �     G
  ��  @      browser_cdl.c str_casecmp get_element_style default_style inline_style add_box_run box_run_count box_runs parse_color.part.0 sys parse_size.part.0 parse_size parse_border_style get_element_type tab_count tabs current_tab url_cursor_blink url_cursor_pos text_run_count text_runs handle_text in_script skip_depth dom_node_count dom_nodes current_element script_buffer_len script_buffer parse_inline_style.part.0 execute_script_content.constprop.0 handle_end_tag handle_start_tag parse_html.constprop.0 parse_state document page_cache link_region_count cache_count history_count history_pos history link_regions navigate.constprop.0 search_mode menus.0 .L19 .L1127 .L1284 .L1287 .L1346 .L56 .L55 .L54 .L53 .L52 .L57 .L50 .L49 .L48 .L47 .L46 .L45 .L44 .L43 .L42 .L41 .L40 .L39 .L38 .L37 .L35 .L36 .L34 .L33 .L32 .L31 .L30 .L29 .L28 .L27 .L26 .L25 .L23 .L22 .L20 .L1095 .L1094 .L1093 .L1092 .L1091 .L1090 .L1088 .L1296 .L1358 .L1357 .L1356 .L1355 .L1354 .L1353 .L1352 .L1351 .L1350 .L1349 .L1347 camel_framework.c initialized.0 temp_menu_count temp_menus js_engine.c str_eq alloc_value next_token keywords operators current_token advance_token eval_binary_op.isra.0 obj_idx.3 static_objects.2 arr_idx.1 static_arrays.0 parse_primary parse_expression parse_statement .L512 .L518 .L517 .L516 .L515 .L513 __x86.get_pc_thunk.si __x86.get_pc_thunk.di _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.dx __x86.get_pc_thunk.bx __x86.get_pc_thunk.bp _GLOBAL_OFFSET_TABLE_ js_console_warn parse_plist_xml js_array_length cm_dialog_input js_new_null js_document_querySelectorAll cm_dialog_render action_count cm_dialog_handle_mouse cm_bind_action nav_home js_new_string js_clear_error js_array_get js_new_boolean js_console_log strncpy_safe fetch_url config_count my_strchr js_to_boolean cm_picker_refresh cm_draw_image current_url cm_dialog_submit cm_dialog_save js_to_number nav_forward cm_init js_get_error parse_menus_from_string js_window_setTimeout on_mouse js_value_ref cm_dialog_open page_offset page_title on_input js_value_unref cm_draw_image_clipped js_new_undefined js_object_set cm_dialog_up_dir cm_get_config js_new_object js_new_array cm_dialog_click actions content_len js_window_alert js_register_native switch_tab js_new_number my_strstr execute_action_by_id cm_load_app_config cm_picker nav_back on_paint js_document_querySelector page_content js_document_getElementById js_array_push cdl_main js_register_dom_api js_get_global js_to_string js_eval js_console_error js_window_setInterval js_set_global cm_dialog_init cm_apply_menus cm_dialog_select_dir my_memcmp js_init open_url_new_tab internal_menu_callback js_object_get status  .symtab .strtab .shstrtab .text .rodata .gnu.hash .data .got .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_rnglists .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                            ��                 !         ��  ��  �                  -         X�  X�  `  
             )   ���o   ��  ��  �  
             3         `�  `�                    9         x�  x�                    >         ��  ��                   G         ��  ��  �                 L         �� �� �                U         ,� ,� 0              ]         \� \� �                 e              � x�                 q              hm �                               �} ;�                 �              + `                  �              � �                 �              I g�                 �      0       �� �                �      0       ��                 �              �� �&                 �   	      �� �� �  
                           �        �         	              �. N
                               �8 �                  