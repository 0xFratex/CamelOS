ELF              �  4   �2     4    (                 @�  @�           Č  �|  �|  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      UWVS����5  ��`>  �t$,�l$0V���!  ���   �É,$���!  ���   ��9�~%�����!  U)��V�Rl����������[^_]�1���[^_]�f�UWVS��4  �K5  ���=  ��4  �l$�E     ��x���P���  �|$$W���!  �PdY^������P��T  �t$(V���!  �PdXZ������P�G P���!  �PdYX������P�F@P���!  �PdXZ������P�G@P���!  �PdY_������P���   P���!  �Pd�E    ��j �l$(U������P���!  �P(�����{  ��1��������D$�������D$�v �E ���I  <.�A  ��U���!  ���   �����%  ���t$�P��T$�D(�P���!  �Pl������   ���t$U���!  �Pl������   ��������PU���!  �Pl������   ��������PU���!  �Pl������   �D$� ��	��   Rj j ���L$$�P���!  �P\���t$U�D$ ��T$���ЋL$$�P���!  �P`YX������P�D$ ��L$���ȋL$(�P���!  �PdXZU�D$ ��T$���L$(�D

P���!  �Pd�D$$� ���v F��@9��������,  [^_]ÐUWVS��   �$ �� ��2  ��z;  h   j ��4   �D$P���!  �P\��j@�l$U���������!  �P(��   �    ����~:���D$�E ��t<.t��H�
���t$�   �ǉ���@�D$9�uύ������8�u������� ������   �     ���!  ���   ���!  ��  [^_]Ív UWVS��\�2  �ä:  �D$x���!  �D$|���!  ���!  ���   ;��!  t�������j���$�   ��$�   ��$�   ��$�   ���!  �P@��h����j(��$�   ��$�   ��$�   ���!  �P@��h����j��$�   ��$�   ��'P��$�   ���!  �P@��$�   �x
��$�   ��
�D$ ��jj�jjWP���!  �PT���!  �PD��x  �� �����  �   ��D$�D$t�hQ������QU�D$|�HQ�ҋ�$�   �p(XZjj�jjWV���!  �RT���!  �RD�� ��t  �	�D$9�7  �   �P��[���PU�D$|��0P��_]jj�j��$�   ��ZP��$�   ��P��$�   ��KP���!  �PT����$�   ��dPh   ���������$�   ��P��$�   ��UP���!  �PH��$�   �h(��h������$�   ��(Ph�   U��$�   ���!  �P@�� h����������P�D$|��2P�t$���!  �PD��$�   �x������D$,�$jj��$�   ��FPW���!  �PP�� h   �������P�D$|��JPV���!  �PD������$jj��$�   ��dPW���!  �PP�� h   ������P�D$|��hPV���!  �PD������$jj��$�   �   PW���!  �PP�� h   ������P�D$|�   PV���!  �PD��$�   ���   �t$8��$�   ��j����|$4�$����jWUV���!  �P@��$�   ���   �L$8�� hfff��� ���P�D$|��.PQ���!  �PD�$����jW��$�   ��?PV���!  �P@��$�   �h@��   �D$$�� � ����  �D$|D$t�D$�|$|W�  �D$p�   �D$��4   1��������D$�������D$������D$ ��4  �D$,�<$�   f��|$��V���!  ���   ����~%��������R�D0�P���!  �Pl����u��������Wjj�EP�t$$���!  �PP�}�� �D$�$9t}h   �VW�t$$���!  �PD���E�$�$�|$9��   ��@��/�T$9���   �ŋD$�$9u��h�׳�j�t$8U�t$D���!  �P@�� �F0�!����|$ ������j�jh�   �EP��$�   �   P���!  �P@�� h   ��t$0W�D$|�   P���!  �PD���L���f���   �����   �������?��=  ��   ��  �l$p*��  �t$t2��jh����Ph�   VU���!  �PT��h����jh�   VU���!  �P@�F�U
�T$ �� �?���  �|$8��t����   �t$8�Ǎl$Pf�h   ��6W�t$���!  �RD������9�uލ�  ����c  �D$x-�   ��������D$p�<��4  �$��	ȍ,�(   �t$|)����������t$tƃ�jh   @Uh�   ��$�   �DP��$�   �DP���!  �PT��jh����Uh�   VW���!  �PT��h����jh�   VW���!  �P@��h����jh�   �D5 PW���!  �P@��h����UjVW���!  �P@��h����UjV���   P���!  �P@�� h   ���A���P�F
P�G
P���!  �PD���$� ��~:�G�D$��$���  1�v h   �WV�t$���!  �RDE���� ���$9(ۃ�\[^_]Ív ����������f�������V���f��P   ����f�h   ���%���RP�|$W���!  �PDh   ���0���P�F PW���!  �PD�� h   ���9���P��:VW���!  �PD������f�UWVS��  ��)  �Á2  �������>���   ��$  �����   ���������|$W���!  �Pd�<$���!  ���   ���|/t$���!  �hd��W���   YZ������R�P�Ճ���W��$  U���!  �Pd���!  �Hd�L$���������T$�<$���   ZY�T$R�P�L$�ы��!  �Pd�T$�,$���   ZY�������P�T$��XZ���!  UW�P4���������  [^_]�f�S����(  ��k1  ��  ���uU�������8�tE�|$
ts�|$tt�|$tI�D$�� ��^w$��$  ����H�
��4  �\$��D ��[Ã|$u��     ��[�f���$  ���~�H���4  � �̐�?����Đ� �����1���붍v VSR�(  �ô0  �D$��x_��   9~U�����������������������P��4  V���!  �Pd�4$���!  ���   ��$  ���   �     ��X[^Ív UWVS��  �'  ��10  ���!  �@d��$�  ���g  ��%�����R�|$<W��Y^�������D$P��$�   V���!  �Pd�4$���!  ���   �����   /t$���!  �hd��V���   YZ������R�P�Ճ����!  �hd��V���   YZW�P�Չ4$���!  �P8������  �D$   �l$(�|$P�������D$�������D$��   ���U�t$��YX������PW���!  �Pd���!  �Pd�T$ �<$���   ZYU�P�T$ �ҋ��!  �Pd�T$ �<$���   ZY������Q�P�T$ �҃����t$V���!  �Pd�4$���!  ���   �����   /t,���!  �Pd�T$��V���   ZY������Q�P�T$ �҃����!  �Pd�T$��V���   ZYW�P�T$ �҉4$���!  �P8����t�D$���!  ���   ��$�  ���������U�t$��XZ�t$ W���!  �Pd���!  �Pd�T$ �<$���   YZU�P�T$ �ҋ��!  �Pd�T$ �<$���   YZ�t$$������v ����$�  V���!  �P,�'����Ĭ  [^_]Í���������S����$  �×-  �D$��u�T$��t%�|$t2��[Ð��u��D$��u��������[Ð��j��������[�f���j ���������[�f�UWVS��  �$  ��%-  ��$0  ���F  ��   9�8  ���!  �H\��4   �����D80�'  Ph   j �t$V��XZ������V���!  �Pd�4$���!  ���   ����~ �|/t��������Q�P���!  �Pd�����!  �Hd�L$����׃�V���   ZYW�P�L$�у���$4  ���x  ��W���!  ���   ����~#��������Q�D�P���!  �Pl������  ��������PW����������u��������PW���������)  �����!  V������R�P����  [^_]Ív Vh   j �t$V��XZ�������D$PV���!  �Pd�4$���!  ���   ����~ �|/t��������Q�P���!  �Pd�����!  �Hd�L$��V���   YZ���S�P�L$�э�x  �����'@���V�������P���!  �Pd���t  �����V�t$���!  �Pd���Y�������  [^_]Ív ��  �    ���������  [^_]Ð��������PW�<��������������������PW�!��������������������PW���������������������PW����������k��������!  V������R�P���f��������!  V�P���Q����v UWVS��  �g!  ��	*  ��$0  ����   ��4  90��   �������} ���   Wh   j �|$W���!  �P\XZ������W���!  �Pd�<$���!  ���   ���|/t,���!  �Pd�T$��W���   ZY������Q�P�T$�҃����!  �Pd�T$�m ���������W���   ZYU�P�T$��]XW�������V���!  �P��  �     ����  [^_]�f�S���]   ���(  ��x  ���~'H����������P���������!  �Pd�9�������[ÐS���   �÷(  ��x  ���t  ;}'@����������P���������!  �Pd���������[Ív UWVS��  ��  ��a(  ��$0  ��  �D$�8����   ��4  �8���!  ���!  ��$8  ��   �?��,�(   �l$���   �������)��������T$����~91����   �,$f�9�| 9$|9�$4  |�j;�$4  �Y  f�@��9�u�9�|���   9�|�t$9�$4  ��  ��D$�     ��  [^_]Ív ��   �����   �������8���  ��$8  ��  ��$4  '~����   ~���$4  ��@x�����*�������)؍�   9�.  ��$8  �+  ��$8  �l���������9��  ��W������$8  �H�����  +�������] ����  ��   ���   ��   ��  ��$4  +
9���   ������*�������)ȃ���%  ���C  ����  ���F  ����   ���������\$S���!  �Pd�$���!  ���   ���|/t+���!  �Pd�$��S���   ZY������Q�P�T$�҃����!  �Pd�$�m ���������S���   ZYU�P�T$�҉$���!  �P0��� �������    �������$4  '��   ���   �M�����$8  �������$4  ��G����  ��$4  ��e����  ��$4  -�   ���������������W���������!  �Pd��x  �����@���W�������P���!  �Pd���t  ����Y������[������$8  ��   ������� �����;����D$�;�$4  �(������������������P   �������$8  ������A�����   ��(��������������������P���>�����������   ������� ������  ���  ��$4  ����!  ���   9�|-�   ����!  ��$4  ��O9��$�����U�
������������Z��������������   ����������������  ���  ��$4  ����!  ���   9�|-�   ����!  ��$4  ���   9������-�   �������������(�����j P�����������������   ����   ��������������x�����j S����������c���������������������P��4  S���!  �Pd�$���!  ���   ��$  ���������jS��������������j���f������������j ���R����������f�WVS��  ��  ��z"  ��$  ���!  h   �t$V�P�4$���!  ���   ����}  ��V������V���!  �Pd����x  �     ��t  �     ��V���������!  �Pd������e���XZ������������������h�  h�  ������P���!  �P<�ǃ���4���P���  V���!  �Pdǃ�     YX��%���P�FP���!  �PdXZ��0���P�F<P���!  �PdYX������P�FlP���!  �PdXZ������P��   P���!  �Pdǃ�      YX������P��  P���!  �PdXZ������P��   P���!  �Pdǃ�!     YX��9���P��  P���!  �Pd������jVW���!  �PX��������   [^_Ã�������P�x����VS�t$��t&�D$�T$��f�@B9�t��8�t���)�[^Ð1�[^Ív UWVS����  ��p   �t$0��tr�L$4��tj���t$<��T>  ���   ��Z�t$@��T>  ���   ��)�x=1��ŉ|$��v F�D$9�'�|$0�PU�t$<W�Q�������uމ����[^_]�f�1���[^_]ËD$�L$��u	�f�9�t
@���u�1�ÐS���  �û  �D$��4:  ��uoǃ4:     ��T>  ����4���R���h@  j ��������T>  �P\���7  �     ���.  �     ǃ8:      ��T>  �������T$ � ��[����t� ��t������T$��[��f���[Ív VSR�z    ���7  ���0����T>  �t$�ҍ��7  ��P�Qd����L$$�L� @���X[^�f�UWVS���  �ø  �D$0�D$���7  ���~N���7  �D$��1��
f�E��$9.~4���t$W��T>  �Pl����u��D� �T$�D� ��t��[^_]���v ��[^_]�S���  ��?  �T$�D$��dt@��etS��x9�8:  ��[�f������ ����D��T:  P�1�������[Ð��������P��������[Ð����	���P��������[ÐVS�L$�t$�\$1����f��@9�t���u��� [^Ð�� [^�UWVS��@��  x  �D$�\$Tǀ8:      h   j ��T:  �|$(W�ǋ�T>  �P\���; �5  ��������|$$������D$(�T:  �D$�f��]�} �  ���t$,S�\$�z����Ń�����  ���t$0P���^�������t��p��8:  ����  �S��8:  �P����  �����D$�1��f�F@�T����t
��"t��u����߉\$ ؋L$� ���\$��"���PU������D$ �����M  9��4�����*����D$߉l$,�f��D$��8�   ���D$9��  ���t$ V�\$�����ƃ�����   9D$��   �D$��8�   ����   ����0���PV�R���������um���\$��8���PV�5����������p����P���e����D- �(���D$ ËD$�1���v ���?���@�T�T���.�����"u��$����P��t��\- ����D$ ËD$�1��@�T�T���b�����"�Y�����u��O����l$,�]�} �������<[^_]�1��n���U��WVS��L�D  ���  �E���.  �M��    �8 ��  ��=����}���[����M����.  �}���E�� �B	�z	 �b  ���u�P���������K  ���u�P����������4  �p����C���PV����������  W��)��~�   �E�RV�}�W�q���Y^��J���R�E�P����������   ���u�P����������   �p����S���PV�j���������   �Eċ ���(����U���W�����M��P��T>  �Pd���U���)�=�   ~��   �U�PV�Eċ �����M��D P�����XZ��]���PW��T>  �Pl�����U���������Eċ �����M��D P�������U�������e�[^_]�UWVS���  ��   ���.  ���~N1�1ۍ��.  �D$�f�C��   9~1���t$8�D$�P��T>  �Pl����u׋D$�D ��[^_]Ív 1���[^_]�f�UWVS��   �  �å  ��$�   ��j���P��T>  ��4$��T>  ��������,$��T>  �_XV�|$W��T>  �Pd�<$��T>  ���   ����~�|�/t��������R�P��T>  �Pd����T>  �pd��W���   ZY������R�P���$   ��T>  �P�ƃ�����   Ph   j V��T>  �P\��h�  VW��T>  �P ����~>� ��V�����4$��T>  �P��T>  �������$����   �Č   [^_]Ð��������P��T>  ��<$��T>  ��,$��T>  ���T>  �4$�P��1��Č   [^_]Ã���T>  ��\���R���1��܍v S���    �L$��T>  ��t#��t��8:  ��~������S��T:  PQ�RX����[�S�D  �  �\$�T$�L$��T>  ��t�@L��t�\$�L$�T$[���[�f�S�  �  �\$�T$�L$��T>  ��t�@L��t�\$�L$�T$[���[�f�UWVS��8�  ��X  ������P��T>  ���T>  ������  ���!  �|$Ǉ�      ��h   �P�ƃ����g  Ph   j V��T>  �P\��j@V�G(P��T>  �P(������  �D$    ��T>  ��\����|$�������|$�t$�T$f��> ��   ���t$V�Pl������   �~0����T>  ��u7���t$�L$���   U�Pl�����  ��T>  �L$���    ��   �L$���  ��?F�i�T$���  ��V�,	����T$���   Q�Pd�T$Չ�$  �F(��(  ����T>  �D$�T$��@9T$�.����t$��V�P�D$ǀ�   ����ǀ�       ��T>  �������$�����,[^_]Ív ��V���   �D$,�,$��T>  ���   ��9D$�y�����U�L$()��P��T>  �Pl�����W�����T>  ��������T>  �_����VS���  ��&  ��T>  ������R�����T>  h   j ���!  V�P\�    ��T>  �������$���[^�f�UWVS���.  ���  �D$ �l$$�|$(���!  �   �C    ��T>  �Rd��tb��P�CP�ҋ�T>  �@d����tX��U�S(R�Ћ�T>  �@d����t6��W���   R�ЋD$<���   ƃ�    ���������[^_]Ð��L���떍������������VSQ�v
  ��  �t$�t$ �t$ �t$�t$�!������!  �@   ����t��T>  �t$�   �D$�BdZ[^��f�X[^�UWVS���
  �Ǹ  ������S���!  �n(U��T>  �Pl����t=��U��T>  ���   ����~-�P��|'/u�E�Ht)�T(��/u��D( ���������[^_]�u�V)�����u���S�F(P��T>  �Pd����f��D' ��1�븐WVS�r	  ��  �����!  �~(W��T>  ���   ����~ �|'/t��������R�P��T>  �Pd����T>  �xd����(V���   ZY�t$�V���D�����[^_ÐUWVS��   ��  �Ƒ  ���!  ���   ��x;��  �  ���C(P�l$U��T>  �Pd�,$��T>  ���   �ǃ����  �|/t6��������R�T$U��T>  �Pl����t���T$R�W��T>  �Pd���{��tb�����   W��T>  ���   ����t7��T>  �pd��U���   ZYW�P�֋��   ����t	��U�Ѓ��    �Ĝ   [^_]Ív ���   ��x�;��  }���T>  �pd��U���   ��XY�?������   P�R�f�� �����$  ������������   P���������f��!�����������PU��T>  �Pd���{�������c����v UWVS��,�J  ���  �|$@�t$D���!  �E ���C  ��T>  ���[  �L$H��p������T$����L$�T$L���������1�T$��jh   @h,  h�  �LQ�L$ �TR�PT��jh����h,  h�  �t$,V�|$$W��T>  �RT��h����jh�  VW��T>  �R@��h����jh�  ��,  RW��T>  �R@��h����h,  jVW��T>  �R@��h����h,  jV���  R��T>  �R@�|$(��
��jh����jj�V
RW��T>  �RT�t$4���� h   �������RV�D$�PR��T>  �RDh   ��URV�D$$�P2R��T>  �RD��h�   hfff��U(RV�D$$���   R��T>  �RH�t$4��(�� �}��  �D$
   ��   ��j�P�D$h|  VW��T>  �R@��h����jh|  VW��T>  �R@��h����jh|  �D$�PW��T>  �R@�D$4��*�� 1�������L$������L$�|$���g�v �L$�D$��jjW�D$�PRQj ������ h   ��D$������   P�GP�D$��#P��T>  �PD�D$�D$�����L$9�td�t$��   9��  ~R9��   u'��h�׳�jhz  �G�P�D$$��P��T>  �P@�� �6�0����$  ���C����L$�>���f��D$��  �}��   �L$�D$���   h   �������RW�t$�VR��T>  �RD�D$$�   �t$��<�$����jh�   P�D$ V��T>  �R@��h   �jh�   �D$PV��T>  �R@�� h   ����   RW�t$�VAR��T>  �RD���L$��jh����jj<Q�L$ �|$$���   R��T>  �RT�t$4��  �� h   ������RV��  R��T>  �RDXZjh�z �jj<�L$Q��@  R��T>  �RT��T>  �RD�� �}t<��L���j�PV�D$O  P�҃��   ��,[^_]�f��D$   ��   �G���f���������1���,[^_]�f���  ��S  ���!  � ��t1���T>  ����Ív UWVS���  ��$  �T$8���!  ���tg�D$0-�  ��9�S���  9�|I�|$4��,  ��;|$<7��,  ;t$<|+�p	9���   �p(9�|)�w	;t$<} �w;t$<|�����f��   ��[^_]Ív �q�t$N�
  ��   ��|  9�|�o(9l$<|v�;t$<|n�T$<)�����������   x�9��  ~�9��   ��   ���   �|$u�k�0��$   �x���PP��T>  ���   R���   R�Pd���V���f���  ���   9�},��6  9�|"9t$<�0�����  ;l$<|�    �������?  9��
���|  9������9t$<�������  ;|$<������������������   �����k�0��$   u�|$ �>����у����   P�4���������S���   ��?	  ���!  ���t�|$tn�|$
t�{t�   ��[Ív ���e�����v ����T>  ���   R���   ���|$t0�L$�Q���^w���>��L$���   Ƅ�    �f��    뗅�~�Ƅ�    뉋$Ë4$Ë<$Ë,$Ë$Ë$�  Terminal /usr/apps/Terminal.app Files /usr/apps/Files.app TextEdit /usr/apps/TextEdit.app /usr/apps /usr/apps/ terminal < FAVORITES Desktop backpack Apps hdd_icon Root Name New Folder New File Refresh Open With: Open Open With... Rename Duplicate Get Info Delete New File.txt New Folder ( ) New File ( ).txt .c .h .md .cfg .json /home/desktop Finder Close Copy View [FW] cm_init: Done.
 fs_new_folder fs_new_file <Menu name=" </Menu> <Item label=" id=" <key> </key> <string> </string> CamelMenuDef [FW] Loading config for:  Info.clist [FW] Picker Refresh...
 [FW] Picker Refresh Done.
 * [FW] Dialog Init...
 [FW] Dialog Init Done.
 /home Save ^ Name: Cancel  [FW] WARNING: cm_init called twice!
    [FW] cm_init: Setting up framework...
  [FW] Failed to allocate config buffer
  [FW] Config not found (or empty):   [FW] Config loaded successfully.
   %   B   '   .       9      )          0             $         1   @                       8   >            <   6      %      -                          !   5   
       (       2   "      #                         ,                                                  3             =       *                 7   ;                /   ?   	   A              :      &       +       4               %         	   Z �J � + �  �@  pB��� � "�(�$W�(B  �   � @  &                                                    !   %   &   (   )   *   -   .           2   3   5   7   8   9   :   ;   ?   A       \O��2�?��� wp�t�k��Lʽ|����h#��*!@�bϐ��Z�-!@������%�CP��"tz5���T*����rMw9J/q|aI�b*�|EI�%`�e�"7{�F?r�v �+R��~c�	�P�Y�^47(2ӏigs�R1�sa��?f��)��͎c* c��Wm+�c%1hjі��=�����"Sn7���K%Gz{1�k�a�M��� �D��	9�xy��Bd8����d�iB���YIE��Q�4                            �6  �6  �6  �6  �6  �6          Files                                      ����������������    /home/desktop                                                                                                                                                                                                                                                   @=  �R  �  �   S  �  `v  �  �N  $   �>  �|                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                89  ���o�:     l�     L}  
   K           ��     �               ���o                                                           	   p   k      �   �    �  `v  @    �  P,  {     >   �>       �  �   8     �   �        3  %       �  j     �   �R       E  @m   	    S   �>       �   �R         ,  �    _   4=       �   �         @Q  @    �  �*  �     @  T      �  �  �     ;  $5  �     �  @v       �  (  3      t.  �    m  �'  :     �   �R         8      #   S   
    �   0=       �   �R       e  �  �       �N       �   �  �     �  �  |     �   `       �  <*  V     �  X  N     �   �R  @     l   8=       Y  �  M     �  �  �     1   �  �     �  �       �  �,  �    �  $   �     /  @%  v     +  ,=       n  �  �    P  L'  D     �  L+  \     =  �%  �    '   �N  �    �   �R       �   �  y     �   �R       P  d  G     +  <3  �    �  �+  �       x#  �    _  �'  :     y   �R       w  �  5     F   @=       �   m              n      has_ext scan_apps app_count app_names app_paths refresh_view entries current_path entry_count renaming_idx selected_idx ctx_active on_paint hist_idx hist_max rename_buf ctx_target_idx ctx_x ctx_y open_with_active commit_rename rename_len on_input start_rename create_item menu_cb open_item history open_with_target_idx launch_with_app nav_back nav_forward on_mouse cdl_main my_memcmp my_strstr my_strchr cm_init actions action_count config_count cm_bind_action execute_action_by_id internal_menu_callback strncpy_safe parse_menus_from_string parse_plist_xml cm_get_config cm_load_app_config cm_apply_menus cm_draw_image cm_draw_image_clipped cm_picker_refresh cm_picker cm_dialog_init cm_dialog_open cm_dialog_save cm_dialog_up_dir cm_dialog_select_dir cm_dialog_submit cm_dialog_render cm_dialog_handle_mouse cm_dialog_click cm_dialog_input  �<     �<     �<     �<     �<     �<     @>     D>     H>     L>     P>     T>     X>     \>     `>     d>     h>            %L             �        2     z   E   &�   	S   X   r   r   r   r   r    'int �   
�   �   �   r    �  �   �   �   r   r   r    \  �   �   �   r   r    0   �      �  #   
    2    �  (  
  ,  2    ) 	^  �   
^   �  4n  �   	r   � 
  n  2    
�   ~  2    �  ,  �	E     U       p    �  �   �  �  �  �    �  *  !�  �  "�  �  %   �  &  $F  '"  (  (;  ,�  )�  0|  *�  4e  +�  8�  .h  <�   /�  @�  0�  D�  1�  H�  2�  LD  3  P�  46  T.  5Z  X�  8t  \0  9�  `�  :�  dZ   ;�  h   <�  l�  =�  p�  >�  t!  ?  x�  @�  |   A-  �  BA  �  CV  ��  F`  ��  G`  �V  H`  �N  I  ��  J`  �u  M  �-   N�  �!  O�  ��  P�  �'  Q�  ��  R  �  S8  �A  T[  �=   Uo  ��  V�  �  W  �k  X  �  [�  � P  P     E  E   i  i     Z  E   �  E   i   u  �  E    �  *�  r   �  P   �  r   �  P  P   �  �  �  r      �  r     P  �  r    �  r   "  P  E   r    	  r   ;  P  r    '  9   h  P  r   r   G   y   �    @  �  r   r   r   r   r    m  �  r   r   P  r    �  �  r   r   P  r   r    �  �  r   r   P   �    r   r   r   r   P   �  6  r   r   r   r   r   r      U  9   U  r   �    ~  ;  t  E   r   i   _  �  E   �  i   �  +y  �  �  P   �  �  �  P  i   �  r   �  P  P  i   �  �  �  P  r    �  �    P  P   �  r   -  �  P  ,   i  A  P   2  V  r   �   F  -&   [  z  z  z  z   r   e  r   �  r   r   r    �  r   �  r   �  r    �  r   �  r   �  i  r   �  r    �  r     r   �  i  r    �  r   8  r   E   i  r   E   z     r   [  r   E   i  r    =  r   o  r    `  r   �  �  �  �   t  m   ]�  $_	�  �   _   �  _'E     �   _3�  ,`		  �   `   �  `)r    7  `6r   $�  `R	  ( �  �  `]�  	  �  
  7	  2   ' 
  G	  2   ? 
  W	  2    sys "	  `  
  w	  2   � 	v  g	  @=  
  �	  2   	2   � 	t  �	   S  	�   r   �R  	4   r   �R  	7  r   8=  	  r   4=  	�   7	  �R  	b   r   �R  	�  r   �R  	  r   �R  	�  r   �R  	(  r   0=  	   r   �R  	  r   ,=  p   &   `  o  #r   `  P  $r    `  
  �
  2   	2    	\  (�
  @Q  
  �
  2   	2   ? 	F  )�
  �N  	�  *r   �N  @,	e  �  -
'	   2  .&   (&  /&   ,�  0e  0.res 1l  1�   2|  4 �  
e  |  2    
&   �  2    9  3  
�  �  2   ? 	�  5�  �>  	�  6r   �>  >  	   =  /  	  �  �  �O  api '"	  � �  
g	  ��}win #E         X	  %O   ]  r    w  �   
~  _  2    !(  
  m 
r   i 
r    "�  ��    ��  x �r   � y �r   �w �!r   �h �(r   �#�  �r   (#  �r   �py �	r   ;      lx �	r   �   �   ly �	r   �   �   V  �	r       k  �  {  i �r   :  2       �P  ^  \  len �r   h  f         cw �r   t  p  ch �r   �  �  cx �r   �  �  cy �r   �  �  �	  ?   �  ��  �H�	  .   k �r   �  �     �	  c  }  bx �r   �  �  bh �r       by �r   $     �  r   9  5    F   i r   P  L    �  �   
P  �  2    "  �  �  ��  x r   � y r   �btn !r   ��  _	r   h  `    `	r   �  �  �  ~	r   �  �  idx �	r   *    n   �  bh r   _  Y  bw r   �  �  bx r   �  �  by  r   	    ~   �  $r   j  b  �   i &r   �  �  �   V  'r   �  �    J      �   �  rx ;r     �  ry <r   �  �  h =r   9  7  �   �  Ar   S  A     �   e  �  Pg	  ��}x  ��}�  ��}�  �   C  �  U  p  �  p  �  h  �  h    �   �  ry lr   �  �  �  mP  �  �  �  �   �  s      �  ,    p   !    key r    0|   �  M   �,  �  �   Q   �d  G   �J  �  �   1f  �p  2�   �r   3f  �
g	   �  �8    �h  idx �r   �  �  �r   �f  �
g	  ��}�   �	r   �  �  �  ��  �  �  len �	r       c   '    �g	  ��}len �r       4  ��}�  �   
  ��}i  �  �  �  �  �  �  �  �  �    �   �  �,  �  �P   �  �r   � �  �
  ��}~  �
g	  ��}�  �	r   #    2   6  �   �7	  ��}M   �  num �G	  ��|c  ��| =   !  num �G	  ��|�  ��|x  ��| �  ��|
  ��| �  u �  u �  �   �  {�  y   �s  idx {r   �  C   m�    ��    �   �  og	  ��{z  og	  ��}a  u �  ��{�  ��{  �  ^�  �   �  �  `�  ��_raw a	r   7  5  8  A   i dr   A  ?    7  ?p   k  ��  �  A�  ��oraw I	r   N  J  J  �  i Jr   a  ]  Y  k  len Lr   w  q     
�  �  2    4D  8r       n   ��   �  8P  � ext 8,P  �`  9	r   �  �    :	r   �  �   $�  �  �   �I  �  � 5�      '   �  �  �  �  s  �  �    $_  �  j   ��  j  � t  �6_  �    X   
�  j  �  �  t  �  �  
  �     h  .  h   7J  T    �W  � 8c  9J  �    �  �   �W  �  �  :c  ��}   ��}2  ��}   �     4L  p      �    /    2     z   E   5�   	S   X   r   r   r   r   r    6int �   
�   �   �   r    �  �   �   �   r   r   r    \  �   �   �   r   r    0   �      �  #   
    2    �  7  
  ,  2     ]  �   
]   �  4m  �   	r   � 
  m  2    
�   }  2    �  ,  �	D     T       o    �  �   �  �  �  �    �  *  !�  �  "�  �  %   �  &  $F  '!  (  (:  ,�  )�  0|  *�  4e  +�  8�  .g  <�   /�  @�  0�  D�  1�  H�  2�  LD  3  P�  45  T.  5Y  X�  8s  \0  9�  `�  :�  dZ   ;�  h   <�  l�  =�  p�  >�  t!  ?  x�  @�  |   A,  �  B@  �  CU  ��  F_  ��  G_  �V  H_  �N  I~  ��  J_  �u  M  �-   N�  �!  O�  ��  P�  �'  Q�  ��  R
  �  S7  �A  TZ  �=   Un  ��  V�  �  W  �k  X  �  [�  � O  O     D  E   h  h     Y  E   �  E   h   t  �  E    �  8�  r   �  O   �  r   �  O  O   �  �  �  r      �  r     O  �  r    �  r   !  O  E   r      r   :  O  r    &  9   g  O  r   r   G   y   �    ?  �  r   r   r   r   r    l  �  r   r   O  r    �  �  r   r   O  r   r    �  �  r   r   O   �    r   r   r   r   O   �  5  r   r   r   r   r   r      T  9   T  r   �    }  :  s  E   r   h   ^  �  E   �  h   �  9x  �  �  O   �  �  �  O  h   �  r   �  O  O  h   �  �  �  O  r    �  �    O  O   �  r   ,  �  O  :   h  @  O   1  U  r   �   E  ;&   Z  y  y  y  y   r   d  r   �  r   r   r    �  r   �  r   �  r    �  r   �  r   �  h  r   �  r    �  r   
  r   �  h  r    �  r   7  r   E   h  r   E   y     r   Z  r   E   h  r    <  r   n  r    _  r   �  �  �  �   s  m   ]�  �  �  T  0-�  �   .�   �  /r   (2  0r   , 
  �  2   '  �	  &   	r    �
  	r   �	  
  l  
�	  (d   
�	  �  !
�	  �X
  $	r   �P  %	r   �[  (�  ��  1�	  �<�  2	r   � 
  �	  2    
  �	  2   ? 
  �	  2    
�  �	  2   ? 	  3�  =�	  6�	  �  �    �  
  �  �  &   >sys �  �|  $2	I
  &id 3  �
  4�    ^	  5)
  
I
  e
  2    �  7U
  `v  f
  8r   @v  
}  �
  2    S	  :�
  �x  -	  ;r   �x   >�
  &key ?  �  @
�
    
  �
  2   � 2
  A�
  
�
    2    �
  C�
  @m  _  Dr    m  ?�	  O `   @  �r   $5  �   ��  key �r   � �  }  len �r        g5  �    �	  fr   <3  �  ��  	o  fr   � 	P  f$r   �mx f/r   �my f7r   �x i	r   >  ,  y j	r   �  �  �  u	r   �  �  �	  v	r   	  	  fy �	r   4	  2	    }  idx zr   @	  <	  �  {r   g	  _	  �4  �  5  �   !�  ^3  i  i�  �  �	  �	   !�  i3  t  j�  �  �	  �	   �3  #   @�  Er   3  %   �  mx E r   � my E(r   �btn E0r   �  s
  �r   t.  �  ��  	�  �r   � 	  �%r   �	o  �0r   �	P  �;r   �x �	r   �	  �	  y �	r   $
  
  �  	r   d
  \
  �	  	r   �
  �
  
  	r   �
  �
  A�  	r   fy 0	r   �
  �
  "�0  �   S  i r   �
  �
  ^  idx r       iy  r   0  $    (O  g  e  �0  ^    !�  �.  H  �v  �  q  o   '�  �.  S  ��  �  �    (�  ��,  �  ��  f  �
�	  ��~len �	r   �  �  =.  �   #�  �P,  {   �#  		  �'O  � len �	r   �  �  B�,  w �,     C�	  �=  )len �r    Dx  �L+  \   ��  �	  �!O  �  �  �  �4O  �  �  	�  �KO  �	  �eO  �cb �~�  �s+  �   #=	  ��*  �   �  	�	  �!O  � 	�  �4O  �	  �KO  �cb �d�  �++     E�
  �<*  V   �(
  [(  3  ��  F@d�  �  e�   2  f&   (�
  g&   ,�  h�	  0*uid i�	  1�  j�	  2*gid k�	  3�   l�  4 GA  m4  	  o	r   �  �  �
  p�      �  f  u	r   =  1    i wr   t  j  '  �  {r   �  �    �r   �  �  2  i  �  �r   �  �  `  �r   �  �   ;)  F   idx �r   �  �      
&   �  2    +�
  H�'  :   �^  (
  H&
  �  �  �   H8O      x HBr   E  ?  y HIr   `  \  dw HPr   �dh HXr   �cx H`r   �cy Hhr   �cw Hpr   � ch Hxr   �$,(  -��  +�  E�'  :   ��  �
  E
  t  p  �   E2O  �  �  x E<r   �  �  y ECr   �  �  	�	  EJr   �	�	  EUr   �,�'  -��  #�
  "L'  D   �  	�
  "E   �  $�
  �r   �%  �  �o  s  �$O  Vh  
�	  ��~)len r   �  
�  V2  	r   P $�	  �O  @%  v   ��  key �'O  � R%  O   i �r   �  �    %(  ��   �  �2  xml �$�  � ptr ��    �  �   �	  ��  ,  "  �  ��  W  Q  �     �  �r   s  m  i �r   �  �  �  ��  �  �  /  ��  �  �      �
  ��  �  �  �  �r     �  R
  ��      �	  ��  c  Y  "#  H   �  k �r   �  �   "�"  L   �  k �r   �  �   c"  �  �"  �  �"  �   "  �   v!  �  �!  �    %s  �x#  �  �j  buf ��  �  �  ptr ��  �  �    �  ��  �  �  @
  ��  �  �  D  ��  �  �  8  �  �@-
  �r   
    �  ��  /  -  �
  ��  =  7    ��  W  S  �
  �r   n  f  �#  �  �#  �  $  �  ?$  j  Q$  �  h$  �  �$  �  �$  j  ,%  �    H�	  ��   8   ��  I�	  ��  �  �  src �+O  �  �  n �4r   #    i �	r   P  J   JM  m�  .�	  m!r   .�  m/r   Kid }O   /l	  c�  |   �2  id c'O  � �   i dr   k  g    %Y  \X  N   �c  �  \!O  � �
  \3�  � /%	  H�  �   ��  api H�  �  {  �  Ir   �x   0�  &�  �     ��  s &O  �  �  c &$r   �  �   $  �  �  �   �X  �	  O  � L	  3O  �T  	r   �  �  �  	r   �  �  8  8   i  r   �  �  g  X    0�  r   �  5   ��  s1 �  � s2 +�  �n =h  �p1 O  �  �  p2 O      �  &   i h        L�  r   �  Mval !r    N�  $   �   �z  1�  � 1�  �2�  C  =  O�  �    �      mg  �  �  �  �  �  �  3�  �   �   w   �  �   �   P#  �+  �   �31  '#  �+   =  �=  21  �  �  ,         I   :;9I8   !I  H }  4 :!;9I�B  'I  '  ! I/  	4 :!;9I?  
I  H }�  4 :!;9I   :;9I  4 :!;9I�B   :!;9I  U    4 :!;9I�B  :;9  4 :!;9I  U  4 :!;9I�B  $ >  .?:!;9!@|   1   1�B  4 :!;9!I   :!;9I    .?:!;9!'@|   :!;9I    :!;9I  !.?:!;9!' !  ".?:!;9!'@|  #4 :!;9!	I  $.1@z  %%  &   '$ >  (& I  ):;9  * '  +&   ,   - 'I  . :;9I8  /.?:;9'I@|  0.?:;9@|  1.?:;9'   2 :;9I  34 :;9I  4.?:;9'I@|  51R�BUXYW  61R�BUXYW  7.1@|  84 1  91R�BXYW  :4 1    I   :;9I8   !I  H }  'I  '  4 :!;9I�B  4 :!;9I�B  	 :!;9I  
I  ! I/   :!;9I  4 :!;9I�B   :;9I  4 :!;9I�B  $ >  U   1�B   :!;9I�B   :!;9I8   :!;9I   :!;9I�B  U   :!;9I  :;9  4 :!;9I?  4 :!;9I  4 :!;9I     :!;9I�B  :;9!	   .?:!;9!'I@|  !1R�BUX!YW  "  #.?:!;9!'@|  $.?:!;9'I@|  %.?:!;9!'@|  & :!;9!
I8!   '1R�BUX!YW  (.?:!;9!@|  )4 :!;9!	I  * :!;9!I8  +.?:!;9!'@z  ,H}�  -I ~  . :!;9I  /.?:!;9!'@  0.?:!;9'I@z  1 1  24 1�B  34 1  4%  5   6$ >  7& I  8 '  9&   :   ; 'I  < :;9I8  =4 :;9I?<  >4 :;9I  ?4 G:;9  @.?:;9'I@z  A4 :;9I  BH }�  C.?:;9   D.?:;9'@  E. ?:;9@|  F:;9  G :;9I  H.?:;9'@z  I :;9I�B  J.?:;9'   K4 :;9I  L.:;9'I   M :;9I  N.1@z  O1R�BXYW  P.1@|   	            �9�9P�9�;W                      ���#F���P����~���#F����#d���P����~���#d����#����P����~���#�����#�����#��       ��V��������      ��U���#(����#(�       ��U��P��U        ��0�������Q����   ��W   ��P    ��������     ��P����~       ��U����:���U         ��V��px���V��vF�  ��0�       ��W��pl�����D�   ��U     ��V��v\�    ��v���vz�    ��0���U       �.�/(��1�3(��3�4(��4�6(�       �.�/���1�3���3�4���4�6��              �.�.�@��.�.S�.�/�@��3�3�@��4�5�@��5�6�@��6�6�@�             �.�/P�3�3P�4�4P�5�5P�5�68=  �6�6P       �,�-w H#(��3�3w H#(��4�4w H#(�      �,�-ȟ�3�3ȟ�4�4ȟ           �,�,r�~2��,�,r 2��,�-`  �2��3�3`  �2��4�4`  �2�         �,�,p w H(2��,�- `  w H(2��3�3 `  w H(2��4�4 `  w H(2�         �,�-R�-�-��}#��3�3��}#��4�4��}#�      �,�-0��-�-P�4�4P      �-�-p H��}#"��-�-pH��}#"��4�4p H��}#"�                   �/�/Q�/�0� �R  ��3�3Q�6�6� �R  ��6�6� �R  ��6�7� �R  ��7�7� �R  ��7�7� �R  ��7�7� �R  �                  �/�/��R  ��/�0��R  ��3�3��R  ��6�6��R  ��6�6��R  ��6�7��R  ��7�7��R  ��7�7��R  ��7�7��R  �   �/�/P                   �/�0P�0�0r 2&q ��6�6P�6�6P�6�6P�6�7r 2&q ��7�7P�7�7P�7�7P      �1�3�(��5�5�(��6�6�(�      �1�20��5�50��6�60�   �#�#P    �$�%W�'�(W   �$�$P   �%�%P    ��1���!��|   ��P  ��0�     ��P��W    ��0���V       ��P��r�����o#�       )2P2KSdjS     8PPdfP     ��� ���    �!�"2��"�"0�    �!�"��"�"1�     �)�*V�*�*�  �
            �/�/P�0�0P                   �+�,P�,�,
� 
�1&��,�,P�,�-
� 
�1&��-�.P�.�.p�}��.�.
� 
�1&��.�.P�.�.
� 
�1&�        �+�+
�
,1&��+�+w 1&��+�,
�
,1&��,�.
�
,1&�    �,�-�
,1&#(��.�.�
,1&#(�      �,�,ȟ�,�,V�.�.ȟ   �-�.V    �,�-	�u D��.�.	�u D�         �,�,
r a  "��,�-R�-�-a  �.�.R    �+�+� 
���+�+P �+�+�
,�             �"�"Q�"�#�H�#�%�D� "��%�*�
�1&� "��*�*�D� "��*�*�
�1&� "�         �"�"R�"�$�T�$�*�
,1&�"��*�*�
,1&�"�         �$�&V�&�*�T#(��*�*V�*�*�T#(�    �$�%ȟ�*�*ȟ    �%�*D��*�*D�         �'�(Q�(�)�L�)�*�T#���*�*�T#��        �%�&0��&�&�D�&�&P�&�(�D     �&�&V�&�(V            �&�&w~��&�&wj��'�'w~��'�'P�'�'���'�'w~�   �&�&Q �!�!�
�� �"�"�
,�         ��P��W�!�!P�!�!W   ��P     ��� ���      ������    ��@���@�         ��P��V���X���X��V             ��P��R���L���L��P��R          ��0����D��R���D��0�       ��w 1���W��W    ��0���0�     ��P���\   ��P   ��Q     ��� ���            �����S�����S���       �����R��R     �����Q     ��� ���            �����S�����S���       �����R��R     �����Q    ��0���S        ��S��S������S           ��U��P��U���\��U       ��P��V��V       ��S��	�x  1���S      ��0���P��0�     ��P���@     ��V�	�	V         ��	V�	�	v{��	�	P�	�V     ��	U�	�U          �	�	P�
�
P�
�
p��
�
q��
�
q p "#��
�q p "#�        �
�
P�
�
p��
�
q��
�
q p "#��
�
q p "#�    �
�
0��
�P    �
�
0��
�
P   ���     ��P��P   ��P     ��P��V   ��P  ��p v ���p v O-( �   ��P       ��V��P��V     ��P��R       ��p v ���r v ���u�v �-( ���r v �-( �           ��� ��Q��� ��Q���            �����V�����V���           �����S�����S���      ��0���P��P    ��0���U       ��� ��� ���      ��� ��P     �����Q     ozPz�W     ��P��U    ��0���V  5�   5�      0�p � �	p � #�*p � �      ��p 0r 8$"�x  "���p 0� 8$"�x  "����0� 8$"�x  "�   ��R���  ��e�           ��P��p���P��P��P��R��P                  �                     �            �         ������ ���� ���� �� � �! ����� �! ��� �  �!�"�"�" �"�"�%�' �,�-�3�3�4�4 �,�-�3�3�4�4 �,�-�4�4 �-�-�4�4 �/�1�3�3�6�7 �/�1�6�7 �1�3�5�5�6�6 �         ���� ������ ������ ��	�	� ���� ���� ���� ���� ���� �!�!�!�" �"�"�"�" �%�&�&�' �+�+�+�+ �+�+�+�+ �,�-�.�.�.�. �/�/�0�0 +    7   �         I   R   	   	   e   1     7���gu<f& .3 f� �0JhK, ��, XY, X�v�	 � 1 fL	�<% �	�	� �; t t J �� � <� <�f�&X��&����&�J�"� r   ������	  �	g<% J	K t : �f X* �� �g+��"��	 �2 �Z*(,./�f � ���� f X0283$	���9 <h �j ���; <g �i ���; <g #	&2�	�	 	g�		�.v@ _�@ y<	K	� � � �U t	g�:�	h<" n < <	�	>�	�@ ��&*	f	�".f �	Y	�	�t=����u $ �  J  �	f	���	u"�	u��	h1���Y�� ��eY$ ;   � �� �. /���� �}JKf* � f	�g �4 �7 I �4 �	LJ��	 ���	 �.	f�g���	fgfV	vwvt: X, �Y"&X(fu$X qX ) t9 fyt�! J, :  ߄g�~�! J fK��)<� ��vK� � f�� �* �- = �* �� ��	 �	x�� � �w�/)� ��)� � �� �2 �5 E �2 �K � �� �uJj	!����)� ��)� � �=Y X���/ J� veU  � X c� ? r� >+�}t� � f�����"� t. t ��A�t ��&� �, � J ��	  # t  �	�<	f�A	M��h	� t+ t �	��	 �;.	 X���= J��	�u$<	i�	�	�; x�8 �	�P �"� �< �9 ��<f	t.<	fK#��  � f�f�Y! �4 �7 L �4 �KR�� ��"<<f��=���	K	=*<	���h��	K	=*<	���&��	�	�"	�	g	h"�X�f�..�> J( 2� J- X; �)    t" J f' J!"�� ��	f$�f �����0	�0  f	�	��f�	���f/%1� �Z�ft1 1� <X������+<=# �? �B S �? �KY�.� ������	�������2 �i/�# �+ =$J����	!�; �1 f  + ,< t1 `X �	&�<�<% �F���� gfg���& J4 u�% �3 % G�u, 	X �g����1�& J4 u.& �4 1 c� �"�����$ � t Z�$ y�&f/F<�&$ �$  ~�$ z }�$  ��$ ,���	h� �	�L1��0YZ0��YYZ������0�	b  �    <   �         �   �   x   x   e   �   @ �  g	 "     	Y.< J& * <1I/;h! ��K�g	  X.! �  	�f � �t& yX5'��	�	K
 s4!./��	h�����f�/I	r. J . J� qJJ@���Y<f&J�K .�g+h�	 t# f  	u u�" J" p X9�i]^ J�r;<X��	sf�<nf	
�D7k� ' �/ # <   J <+ J/=  	-.=  )7 ���x'��	!<P	��X	/	�	�u>!f�(�11<-h8) - 1I1. J1 X['<�<K��fN�-�<h�"/ ��Ju�!{Y�: $ : < � : t�CG : I$ : J* � �w< $ < < �K?C < I$ < J+ �< � �	J<P2�Y�!�tg�#%1�
�	[<S	�	�	�#	�  �1 	>!	�	�K	��.	�	�#	� �0 	?!	!	�<.�1J��y<z�2. i .�A<  ,;�!	 �# �  	�&tf �7 t> �Js/5��. �K �� f. tv� ��!�"/{L��f��	s�;  S �	�	fgx<.	l�<	f�'�!	f JKf	KL\Xgf J <  J J JK  = |=gf J <  J J JK  = <!�	f�@)��"L	 ���	t<	� �	�2	zd<0 J�= b  �Y,�/J.K+�)� cf J J !v��f�j���g�?Jf< � � � ff�f�<fgf�h���u� J�� t�� t��!uu z� � ���!K� t  f J �= ;KL!	 �s�- � <9 �   + . J
Z%Zu }+ .g J t	�&	Y &-.0<�� t9 t ��)� ��Y�L�' J�K �/ t J, <	u��	| Xu%� � yf/f% t�
f	s�f+ J�%� �h. �	m�8��M<t�t	g��<B��� � f��|��|�	 �.��|��|�	 �.x�M'����J�J$�&	u	I[����
 �E . � J	�w:�	�) pX J J <	�	�	���@X�	@2E� � �	�	���#��('*"� � f���0 O� .�+ ��� .5��� J�;OY�L�{��{�.��{� J fH�{�." �6 f, fi< � <( J" <: f0 <	gYF );XN�t	s[$  f	F( @G f8 .	gfX	[f .��*iS t4 <�.Vft��	if2 J f7 JO �C f	g	gjf1 � X6 �N �B f9 c� �0 s
�0<��E<tf'���LyyxfX	p�u	]<f	��t, XY-�-�	p	g. J: 
 malloc print strcmp sprintf open_with_active socket hist_max close commit_rename nav_back strncpy rename_len kernel_api_t win_handle_t cdl_symbol_t lib_name paint_cb_t input_cb_t free plen app_idx rename_buf exec item_count draw_rect hist_idx dates candidate fs_create on_mouse cdl_main recvfrom menu_cb memcpy scan_apps recv fs_list get_kbd_state menu_cb_t launch_with_app current_path draw_text_clipped entry_count toolbar_h create_item get_launch_args strcpy open_item temp attr force_dialog net_get_interface_info elen strlen process_events bind start_block size selected_idx draw_image_scaled row_y app_names full_path last_fs_gen fs_rename label old_full symbols action_id cdl_exports_t base version ctx_active entries filename get_fs_generation fs_write send start_rename sidebar_w open_with_target_idx exec_with_args direntry_t has_ext GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection http_get history nav_forward list_y unsigned char is_dir fname strncmp counter draw_rect_rounded create_window app_count draw_text exit mouse_cb_t connect icon uint32_t itoa newp on_input sendto set_window_menu exports app_paths win_h mem_total flen fs_exists win_w ping new_full memset func_ptr get_ticks memmove fs_read refresh_view ctx_y dpath list_start_y mem_used menu_def_t target fs_delete on_paint renaming_idx ctx_x realloc dns_resolve ctx_target_idx symbol_count key_content_end hlen cm_bind_action clist_path parse_plist_xml file_buf my_memcmp my_strchr cm_dialog_select_dir file_picker_cb_t perm visible_items start_dir long long int cm_dialog_submit show long long unsigned int my_strstr parse_menus_from_string cm_dialog_input selected_index config_count current_dir cm_dialog_save val_tag name_ptr value initialized real_idx nlen default_name menu_end key_tag short unsigned int i_idx cm_dialog_handle_mouse dirname max_read file_picker_t cm_init temp_menu_count cm_dialog_open needle temp_menus action_bind_t execute_action_by_id strncpy_safe cm_dialog_click title id_p req_h haystack dest menu_idx cm_picker menu_tag req_w cm_dialog_up_dir cm_get_config list_h cm_picker_refresh item_h short int buff klen config_pair_t key_content_start lbl_p scroll_offset action_count cm_dialog_render cm_dialog_init cm_apply_menus func mode val_content_start vlen cm_load_app_config item_tag cm_draw_image_clipped buffer win_handle win_y filter filter_ext val_content_end item_ptr key_name raw_entry_t internal_menu_callback filename_input app_bundle_path win_x cm_draw_image item_idx actions safe_div2 usr/apps/files_cdl.c /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/apps usr/apps/../../sys cdl_defs.h usr/lib/camel_framework.c usr/lib usr/lib/../../sys camel_framework.h     ���� |�  `           n   A�A�A�A�C,T0` G(G,E0F K
A�A�A�A�AEA�A�A�A�  4      p   k  A�A�A�A�F�c�K�J�A�G�K�J�A�G�D�J�A�G�D�J�A�G�D�J�A�G�G�S�B�E�G�L�y�A�O�L�D�L�L�K�D�A�L�K�G�A�L�K�G�A�L�X�B�B�J�L�D�A�V�J�A�G�V�J�A�A�V�R�UA�A�A�A� \       �  �   A�A�A�A�F� G� P� B� K� L� B� E� F� X� yA�A�A�A�t      �    A�A�A�A�Cp{|B�G�G�G�G�L|E�B�G�G�G�L|E�B�G�K�G�dxB|B�B�B�A�A�[p[tGxA|H�M|AxB|B�B�B�A�A�UpZtGxA|H�C|AxB|B�B�K�K�K�L|K�E�F�K�K�V|E�K�E�A�G�LpEtGxH|D�b�B�K�A�LpEtGxH|A�T�B�K�A�LpEtGxH|A�T�B�M�A�LpEtGxJ|A�t�A�A�A�]pEtGxH|A�R�A�K�A�`po|A�OpHxG|E�LpM|A�B�B�D�D�OpPtAxA|D�Lpw|E�B�D�A�D�LpV|B�B�E�D�M�LpEtDxA|J�LpFxB|E�A�E�A�A�L|E�B�E�A�A�VpktBxA|D�Rp^xB|E�A�E�L�L�LxB|E�A�E�A�A�L|E�B�E�A�A�L|E�B�E�E�A�L|E�A�B�A�A�L|E�A�B�A�G�LpEtGxD|D�LpctAxA|D�SpJ
A�A�A�A�DitGxA|E�N�G�D�A�LpEtGxD|A�Lp  �       �    A�A�A�A�F�m�F�E�[�S�A�G�A�G�C�E�C�A�H�o�A�E�C�]�A�F�C�G�A�G�A�F�LA�A�A�A� ,       �  �   A�Cj
A�AP
A�C   0       �  y   A�A�ApJG qAA�A�l      ,  �  A�A�A�A�F�l�A�E�C�A�K�H�[�V�A�G�A�G�C�E�L�A�G�A�A�C�Q�u�A�D�C�A�G�A�`�A�A�C�]�A�G�C�I�C�D�A�[�Z�A�G�A�G�C�I�P�A�G�A�A�C�U�f
�A�D�C�A�D�A�`�A�A�C�]�A�D�HC�G�A�TA�A�A�A�A�����  L       �  j   A�Ce
A�BU
A�BCB HC
A�CCB HCA� �      8    A�A�A�A�F�H�E�B�E�C�A�F�A�[�N�G�C�L�W�A�G�A�A�C�I�R�A�O�H�G�E�L�K�G�A�J�G�G�A�H�K�G�G�F�F
A�A�A�A�DA�E�B�E�C�A�K�A�[�N�G�C�L�P�A�G�A�F�C�Q�K�A�J�V�C�A�D�S�F
A�A�A�A�DZ
A�A�A�A�BC�G�A�H�K�G�A�H�K�G�A�H�K�G�A�H�K�G�G�F�H�G�F� �       T    A�A�A�A�F�y�E�B�E�J�A�F�A�[�W�A�G�A�G�C�I�\�A�G�A�A�C�G�A�A�J�X�FA�A�A�A� (       d  G   A�C]JF QCA� (       �  M   A�CcJF QCA�       �  �  A�A�A�A�F��
A�A�A�A�D/�F�E�[�V�A�G�A�G�C�I�[�A�G�A�A�C�\�y�A�F�T�K�A�J�]���A�J���B�A�J�n�B�A�J�P�L�G�e�H�B�A�J�H�B�J�H�B�J�      �  �  A�A�A�F�]�E�T�K�A�G�L�[�A�F�T�A�F�F�F�E�E�G�N�G�G�T�A�G�D�J�A�G�D�J�A�G�D�J�A�G�G�T�A�G�G�J�A�G�G�T�A�G�G�O�B�A�A�UA�A�A�A����C�G�       �5            �5            �5            �5        ���� |�  ,   �  �  5   A�A�k
�A�BC�A�   l   �  �  �   A�A�A�A�C0^<D@O<D@O0a4A8D<A@H0K
A�A�A�A�CGA�A�A�A�     �  �     D   �  �  �   A�ClG EEBF @A�B�W
A�DCA�0   �  X  N   A�A�AZJM VAA�A�X   �  �  |   A�A�A�A�C0|8D<A@L0W
A�A�A�A�ECA�A�A�A�T   �  $   �   A�Cl
A�CCW HC
A�BCG HC
A�BCG HCA�,   �  �   8   A�A�k
�A�BF�A�   �   �  �   �  A�A�A�A�CTaXB\K`NP}XD\A`NPKXD\A`JPgXK\A`LPAXD\A`NPiXG\A`JPGXK\A`JP�
A�A�A�A�A(   �  x#  �  A�BF�����A�A�A�X   �  @%  v   A�A�A�A�C0w8D<G@L0O
A�A�A�A�DEA�A�A�A��   �  �%  �  A�A�A�A�F�Y�e�A�A�E�Z�N�G�C�K�L�A�G�A�G�C�W�I�E�B�A�L�E�A�A�L�K�A�e�K
A�A�A�A�BC�G�m�H
A�A�A�A�AC�M�E�,   �  L'  D   A�ClAGA FCA�     �  �'  :   A�t
�CA�   �  �'  :   A�t
�CA��   �  (  3  A�A�A�A�CLRPQ@_LEPH@IDEHBLAPLDBHALDPN@@HDLAPF@]HDLKPF@~HALTP[@bLAPo@C
A�A�A�A�DCLAP\@MHALJPL@  4   �  <*  V   A�A�CX EKBG ]A�A� d   �  �*  �   A�A�A�A�C z(A,D0N G(A,D0N G(A,G0]A�A�A�A�B ����  D   �  L+  \   A�A�ASDDD U[
A�A�DAA�A�   X   �  �+  �   A�A�A�A�C(R,J0L G,A0O m
A�A�A�A�AO(A,D0L  T   �  P,  {   A�A�A�NJ ONGC LLD GADC JA�A�A�   �   �  �,  �  A�A�A�A�F�j�D�E�]�R�G�E�L�G�E�C�L�J�G�O�P�A�G�A�A�C�K�G�A�E�L
A�A�A�A�D^
�A�I�A�P�C�DZ�H�J�M�G�A�L�     �  t.  �  A�A�A�A�C@`HBLEPETEXE\I`FHBLEPETEXE\E`LLEPBTEXA\A`LLEPBTEXG\A`LLEPETBXA\A`LLEPETBXA\G`SHBLEPBTBXD\A`S@EDGHALHPNTDXA\H`LLEPETDXA\K`S@ZLBPATIXA\A`LLEPBTEXA\A`LLEPBTEXG\A`S@lHBLBPATHXA\B`H@EDQHDLHPW@eLEPBTEXD\H`L@JDGHALHPbTEXA\E`LLEPBTEXE\A`L@EDGHALHPL@GHBLEPBTBXA\O`V@EDGHALGPJLAHBLEPBTBXE\G`U@NDAHALJPE@H
A�A�A�A�CaA�A�A�A�   �  3  %   T   �  <3  �  A�A�A�A�C0�
A�A�A�A�Dy4A8N<G@F0�<H@H0(   �  $5  �   A�Cs
A�DOM I    �  �5        �  �5        �  �5        �  �5        �  �5                                 ��   `          `          `       #    `       )    ]       1    =  ,     9            ��   �|       K   �x       Y   �x       i   �x                    ��t   �5        �   �5        �   �|       	 �   �5        �   �5        �   �5        �   �5          l>          x#  �    '  @Q  @    1  $5  �     A  �R       G  �  �     T  @=       a  t.  �    r  @v         3  %     �      n     �  X  N     �  �R       �  �   8     �   m       �  �       �  �R  @     �  (  3    �  �'  :       �,  �      L+  \     -  �  j     5  p   k    ?  �R       H  �  M     T  �  �     \  �   �    t  �R       }  �  �    �  �*  �     �  ,  �    �   S   
    �  �R       �  �  �     �  �'  :     �  T      �  0=       �  �+  �       @%  v       <3  �    !  �R       ,  `v  @    4  �  y     A  4=       N  �  �     X  �  |     m  �%  �    �  �R       �   `       �  d  G     �  ,=       �  �      u  @m   	    �  �N       �  �>       �  �N  �    �  �  �    �  �      �  <*  V     �  L'  D       P,  {     !  8=       .  �  5     8  $   �     O  �>       W  8       files_cdl.c sys last_fs_gen win_w win_h menus.0 exports camel_framework.c initialized.0 temp_menu_count temp_menus __x86.get_pc_thunk.si __x86.get_pc_thunk.di _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.dx __x86.get_pc_thunk.bx __x86.get_pc_thunk.bp _GLOBAL_OFFSET_TABLE_ parse_plist_xml app_names cm_dialog_input ctx_y refresh_view current_path cm_dialog_render action_count cm_dialog_handle_mouse has_ext cm_bind_action open_with_active strncpy_safe config_count my_strchr rename_buf cm_picker_refresh cm_draw_image cm_dialog_submit cm_dialog_save menu_cb scan_apps hist_idx nav_forward cm_init parse_menus_from_string hist_max on_mouse cm_dialog_open create_item history ctx_active on_input cm_draw_image_clipped launch_with_app ctx_target_idx cm_dialog_up_dir cm_get_config cm_dialog_click rename_len actions start_rename renaming_idx my_strstr execute_action_by_id cm_load_app_config ctx_x cm_picker nav_back open_with_target_idx on_paint app_count entry_count app_paths cdl_main commit_rename cm_dialog_init cm_apply_menus cm_dialog_select_dir selected_idx my_memcmp internal_menu_callback entries open_item  .symtab .strtab .shstrtab .text .rodata .gnu.hash .data .got .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_rnglists .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                         �5                 !      2   �5  �E  R                -         89  8I  �  
             )   ���o   �:  �J  �  
             3         �<  �L  `                  9         @>  @N  ,                 >         l>  lN                   G         �>  xN  D>                  L         �|  Č  �                U         L}  L�                 ]         l�  l�  K                 e              @�  �/                 q              �  �                               ��  �                 �              ��  @                  �              ��  �                 �              ��  �                  �      0       _ �                �      0        �                 �              � 0                 �   	      ��  ��  �   
                           �' p              	              h- a                               �1 �                  