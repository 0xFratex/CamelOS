ELF                  4   �%      4    (                 4  4           8  8  8  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      1�Ð�2     ��   ��t� f�Ív �     �T$��   ��x���Ë$�                                                      00���M֋                kernel                                �                       get_ticks                           log                                8                        @   ���od            �  
                                   ���o                                                                                               k_get_ticks k_log cdl_main �            $     �	       {             ;       �  1   
0  �   C   �   	P   U   o   o   o   o   o    int �  
�   �   �   o    h  �   �   �   o   o   o    k  �   �   �   o   o    	0�   �  �    �  #       1    
-      #  1     	R  �  
R     4b  �  	o   �   b  1    �   r  1    �   #  	�	  u     �  -  �  F  S  V  �  \  �   p  �  !�  �  "�  �  %�     &�  $:  '�  (�   (�  ,T   )p  0�  *�  4L  +p  8  .%  <a  /I  @8   0h  D�  1�  H�  2�  L�  3�  P�   4�  T(   5  X�  81  \�  9Q  `  :f  ds  ;�  hL  <�  l�  =�  pM   >�  tp   ?�  x   @Q  |2  A�  ��   B�  �  C  ��  F  �C  G  �B  H  �{  I<  �^   J  �  M�  ��  NZ  ��   Ox  ��  Px  ��   Q�  �(  R�  �X  S�  �c  T  �=  U,  �    VJ  ��   W�  �w   X�  �  [\  �          C   &  &   
+    C   F  C   &   2  V  C    K  [  o   p     a  o   �       u  �  �  o      �  o   �    �  o    �  o   �    C   o    �  o   �    o    �  8   %    o   o   E   v   �    �  I  o   o   o   o   o    *  h  o   o     o    N  �  o   o     o   o    m  �  o   o      �  �  o   o   o   o      �  �  o   o   o   o   o   o    �    8     o   �    r  �  1  C   o   &     K  C   K  &   P  6  f  �     V  �  �    &   k  o   �      &   �  �  �    o    �  �  �       �  o   �  �     �  &  �     �    o   �     &     7  7  7  7   o   "  o   Z  o   o   o    A  o   x  o   K  o    _  o   �  o   K  &  o   K  o    }  o   �  o   K  &  o    �  o   �  o   C   &  o   C   7   �  o     o   C   &  o    �  o   ,  o      o   J  �  �  �   1  �   ]}  	$_	{  �  _   �   _'C     V  _3Z  	,`	�  �  `     `)o    �   `6o   $#  `R�  ( {    `]�  �  O  sys �  4  {  �  1       	�  �   B   �  �      �         �F	  api '�  �  �        �y	  msg   �    � �   �  o          �  I   :!;9I8   !I  'I  '   :!;9I  I  ! I/  	:!;9  
$ >  4 :!;9I   :!;9I  %     $ >  & I  :;9   '  &       'I  4 :;9I  .?:;9'I@z  .?:;9'@z  H}�  I ~  . ?:;9I@z                    ;           �     7   �         H   P         b        K�"!f' J8J,J�	� g net_get_interface_info memmove cdl_main set_window_menu draw_text my_exports strchr fs_delete get_fs_generation strstr http_get draw_rect_rounded fs_create win_handle_t kernel_api_t symbol_count sendto func_ptr paint_cb_t menu_def_t dns_resolve strlen bind itoa cdl_exports_t ping strcpy my_symbols long unsigned int close mem_used fs_exists cdl_symbol_t recv mouse_cb_t strncpy get_kbd_state memset exec_with_args draw_image k_get_ticks realloc input_cb_t draw_text_clipped exec action_id get_launch_args item_count process_events items create_window send char sprintf fs_list mem_total strcmp free recvfrom draw_rect menu_cb_t print GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection memcpy exit k_log socket uint32_t fs_rename lib_name fs_read label strncmp draw_image_scaled malloc connect version fs_write usr/lib/syskernel.c /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/lib usr/lib/../../sys cdl_defs.h    ���� |�                                                  ;                                  ��   4          �   ,        �   H                  ��'   8        0   ;         F   (        \           b            k             syskernel.c sys my_exports my_symbols _DYNAMIC __x86.get_pc_thunk.ax _GLOBAL_OFFSET_TABLE_ k_log cdl_main k_get_ticks  .symtab .strtab .shstrtab .text .gnu.hash .data .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_aranges .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                            ?                  %         @   @  $                !   ���o   d   d  ,                +         �   �  �                   1         (  (                   :         4  4                    ?         8  8  �   	             H         �  �  @   	            P                                 X              4  �	                 d              �  c                 r              '                     �              G  �                  �      0       �                  �      0       �"  m                 �              `#  T                  �   	                                        �#  �      	         	              t$  w                                �$  �                  