ELF              �  4   ��      4    (                  0   0            @   0   0  �%  �%           _  O  O  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      VSS�f)  ��0  �t$��8  ��tz��4  ��tpQh �  j R�P\��h��  ��4  V��8  �P ����xE��0  ��4  � ��V��`���P��8  �Pdǃ(      ǃ$      ǃ,      ��X[^�f�VSP��(  ��|/  �t$��8  ��tE��V�P8����t>R��0  ��4  V��8  �P$YXV��`���P��8  �Pdǃ,      ��X[^Ív ��j V��8  �P,���UWVS��  �G(  ���.  ��8  ���  ��$8  ��T�����$<  ��P�����h����j(��$L  ��$L  ��$L  �P@��h����j��$L  ��$L  ��'P��$L  ��8  �P@��$P  ��
�D$0��$T  �z��jj�jj<WP��8  �PT��$T  �p�� h   �������PV��$<  ��P��8  �PD]Xjj�jj<W��$L  ��PP��8  �PT�� h   �������PV��$<  ��bP��8  �PDXZjj�jj<W��$L  �   P��8  �PT�� h   �������PV��$<  �   P��8  �PDY_��`���P�|$|W��8  �Pd����,  ����  hUUU�WV��$<  �   P��8  �PD��$D  ��(�D$$��$L  ��@�$����Q�L$��$L  P��$L  ��8  �P@��$  ��4  �� ���L$�S  ��0  ���E  �
   )�1��D$�����D$�����
   �T$0�T$��$8  ���~   9����
   ����   ��xT9�}P<~L�T$�L$�D$0�D$1 ����$D  h   ��t$ �D$,�P��$L  �P��8  �PH�� �T$�L$�v ��F9�0  |4��4  9�(  u�l$�|$�0<
�g������
   F9�0  }�f���8  �~@�l$���tZ�D$��xR9�}N��   A��   �gfff��������)Ȩt,��h�z �j
j�D$�L$,�P��$L  �P�׃� ��8  ��$<  ��$4  �<��h����j��$L  ��$L  ��$T  �D�P��$L  �V@���t$,V��0  ��8  ���   XZ������P�l$U��8  �PdYXV�D$DP��8  �PdhDDD�U��W�t$,��8  �PD�� ��$<  ��$<  ��$<  ��$<  ��  ����  [^_]�f���8  �hd��W���   ZY������R�P�Ճ��<����v ��8  �D$0�D$������UWVSR��#  �*  �l$��4  ��tZ��0  �$=��  J��(  9�~��>�v �X��H9�u���>G��(  �$C��0  � ǂ,     ǂL�������X[^_]�f�UWVS�U#  ��*  ��4  ��tM��(  ��~C��0  9�}�/�7���X�@9�u��]���(  N��0  �7 ǂ,     ǂL�������[^_]ÐWVS��"  � )  ��4  ��tH��(  ��0  9�}8�q�9�}��L��v �X�@9�u���0  �7 ǂ,     ǂL�������[^_�UWVS�"  ;)  �\$��~x��0  ��4  ��T�����1��
   �
   ��v ��@9�t9�~�| 
t59����   @9�u�\$��t�D$��D$��t�D$�[^_]Ív ���
   뱹
   �
   ��f�UWVS����!  �(  ��0  ����   ��4  ��T������$�T$1���� �
   �
   �|f9�~�<
tP9$~'��@9�|,9\$ u�9L$}/��+t$9�}Ӊ��D$�ː���   @9�}ԋD$��[^_]Ív �t$)��σ��
   �f����� ~Յ��   H�D$�D$��[^_]ÉT$�WVS���!  ���'  �D$P�D$P��(  �f�����P����t$��$  ��)�����	�F���$  �
   �z�9���T��)Љ�$  ��y
ǃ$      ��[^_Ív U��VS���   ��G'  �u�E�P�E�P��(  �������L��������u	�U���L������6��M����
}�
   PR�M�����(  �������e�[^]�UWVS���&   ���&  ��(  �l$0����   ��0  9�~{F�t$��(  9�~l��4  �T$1�L$����
tB�   9���   �Њ�� u�L$�����   ��(  9�~$1���v @�9���   ���< t��t��(  ǇL����������V�����[^_]�f���~�N��(  t؋�4  ��1���v �   Ht<�< t����tJ��(  1��<
t�   Jt�ӊD�< u����t���(  �Ǉ(      �v�����D$�H����v ���UWVS��(��  �Ð%  �t$<V�   ������   ����   �D$    �D$    �D$    ��8  ����   ���   ����   Q�T$R�T$R�T$R�Ѓ����   o����   �F���	��  ���\�����ዃ(  ��0  9�}0��4  1��f�@�   9���  �ǀ<
u����t��(  f�ǃL��������������[^_]Ð���   ��~�F���	��  �����������	��  ��
t6���a  �P����f����   ���~ӍF���	�?  �����������j
������뀐��(  ���b�����4  1���H�C  �ŀ|�
u���>�����(  �3����v �
   �v ��j������Nu��"����v �
   �v ��j��f�����Nu������v ����������f���j�B����������f���j��.�����������T$��t.��j������������D$��t0��j�n���������f���(  ���z���H��(  �n���f���(  ;�0  �Z���@��(  �N���f��F���^�O�����V�_������>����v ��j �J����$    �>���������f�ǃ(      ������S����  �ï"  ������������P������P������P�  ��[�VS����  ��z"  ������P��`���V��8  �Pl����tR��V��8  �P8����t*R��0  ��4  V��8  �P$ǃ,      ��X[^�f���j V��8  �P,���������������P�����P������P�����P�  �� X[^Ív ���  �!  ǀ0      ��4  � ǀ(      ǀ,      ��8  ������Q��`���P�Rd��ÐWVS��  ��x!  �|$�t$��(w)�|$��   ��P���VWP��T�����  ��[^_Ív ��P���~��P�9�~ك|$u҃���$  �Lظ���*�������)ȍ Ѝ�
   PW�N�����(  ǃL���������P�����뇍v �G���<v$�G���<v(��j�����<�_����0����l����v ������_���f�������S���f�S����  �Ë   �D$�T$��u��t��t0��u�������[Ð������[�f���u鋃8  �@��[�������ӐWVS��  �x  ��*   ��$  ��8  h �  �V��4  ����tQh �  j P��8  �P\����V�  �  XZh   �t$V��8  �P�4$��8  ���   �����   ��������������������h�  hX  �����P��8  �P<�ǃ�������P��    V��8  �Pdǃ     XZ������P�FP��8  �PdYX������P�F<P��8  �PdXZ������P�FlP��8  �PdYX��$���P���   P��8  �Pd������jVW��8  �PX�� �����   [^_�f���V����������VS�t$��t&�D$�T$��f�@B9�t��8�t���)�[^Ð1�[^Ív UWVS����  �È  �t$0��tr�L$4��tj���t$<���  ���   ��Z�t$@���  ���   ��)�x=1��ŉ|$��v F�D$9�'�|$0�PU�t$<W�Q�������uމ����[^_]�f�1���[^_]ËD$�L$��u	�f�9�t
@���u�1�ÐS���!  ���  �D$���  ��uoǃ�     ���  ����p���R���h@  j ���������  �P\��`  �     ��@  �     ǃ�      ���  ��)����T$ � ��[����t� ��t��H����T$��[��f���[Ív VSR�j  $  ��`  ���0�����  �t$�ҍ��  ��P�Qd����L$$�L� @���X[^�f�UWVS���  ���  �D$0�D$��`  ���~N���  �D$��1��
f�E��$9.~4���t$W���  �Pl����u��D� �T$�D� ��t��[^_]���v ��[^_]�S���  ��W  �T$�D$��dt@��etS��x9��  ��[�f������ ����D���  P�1�������[Ð����>���P��������[Ð����L���P��������[ÐVS�L$�t$�\$1����f��@9�t���u��� [^Ð�� [^�UWVS��@��  �  �D$�\$Tǀ�      h   j ���  �|$(W�ǋ��  �P\���; �5  ����X����|$$��^����D$(��  �D$�f��]�} �  ���t$,S�\$�z����Ń�����  ���t$0P���^�������t��p���  ����  �S���  �P����  �����D$�1��f�F@�T����t
��"t��u����߉\$ ؋L$� ���\$��e���PU������D$ �����M  9��4�����m����D$߉l$,�f��D$��8�   ���D$9��  ���t$ V�\$�����ƃ�����   9D$��   �D$��8�   ����   ����s���PV�R���������um���\$��{���PV�5����������p����P���e����D- �(���D$ ËD$�1���v ���?���@�T�T���.�����"u��$����P��t��\- ����D$ ËD$�1��@�T�T���b�����"�Y�����u��O����l$,�]�} �������<[^_]�1��n���U��WVS��L�L  ���  �E��@  �M��    �8 ��  �������}��������M���`  �}���E�� �B	�z	 �b  ���u�P���������K  ���u�P����������4  �p��������PV����������  W��)��~�   �E�RV�}�W�q���Y^������R�E�P����������   ���u�P����������   �p��������PV�j���������   �Eċ ���(����U���W�����M��P���  �Pd���U���)�=�   ~��   �U�PV�Eċ �����M��D P�����XZ������PW���  �Pl�����U���������Eċ �����M��D P�������U�������e�[^_]�UWVS���  ��8  ��@  ���~N1�1ۍ�`  �D$�f�C��   9~1���t$8�D$�P���  �Pl����u׋D$�D ��[^_]Ív 1���[^_]�f�UWVS��   �  �ý  ��$�   ������P���  ��4$���  ��������,$���  �_XV�|$W���  �Pd�<$���  ���   ����~�|�/t��������R�P���  �Pd�����  �pd��W���   ZY������R�P���$   ���  �P�ƃ�����   Ph   j V���  �P\��h�  VW���  �P ����~>� ��V�����4$���  �P���  �������$����   �Č   [^_]Ð��������P���  ��<$���  ��,$���  ����  �4$�P��1��Č   [^_]Ã����  ������R���1��܍v S���u  /  �L$���  ��t#��t���  ��~������S���  PQ�RX����[�S�4  �  �\$�T$�L$���  ��t�@L��t�\$�L$�T$[���[�f�S��  �  �\$�T$�L$���  ��t�@L��t�\$�L$�T$[���[�f�UWVS��8�  ��p  ������P���  ����  ������  ��@  �|$Ǉ�      ��h   �P�ƃ����g  Ph   j V���  �P\��j@V�G(P���  �P(������  �D$    ���  ������|$�������|$�t$�T$f��> ��   ���t$V�Pl������   �~0�����  ��u7���t$�L$���   U�Pl�����  ���  �L$���    ��   �L$���  ��?F�i�T$���  ��V�,	����T$���   Q�Pd�T$Չ�$  �F(��(  �����  �D$�T$��@9T$�.����t$��V�P�D$ǀ�   ����ǀ�       ���  �������$�����,[^_]Ív ��V���   �D$,�,$���  ���   ��9D$�y�����U�L$()��P���  �Pl�����W������  ���������  �_����VS���  ��>  ���  ��	���R������  h   j ��@  V�P\�    ���  ������$���[^�f�UWVS���:  ���  �D$ �l$$�|$(��@  �   �C    ���  �Rd��tb��P�CP�ҋ��  �@d����tX��U�S(R�Ћ��  �@d����t6��W���   R�ЋD$<���   ƃ�    ���������[^_]Ð������떍������������VSQ�~
  ��0  �t$�t$ �t$ �t$�t$�!�����@  �@   ����t���  �t$�   �D$�BdZ[^��f�X[^�UWVS���"
  ���  ������S��@  �n(U���  �Pl����t=��U���  ���   ����~-�P��|'/u�E�Ht)�T(��/u��D( ���������[^_]�u�V)�����u���S�F(P���  �Pd����f��D' ��1�븐WVS�z	  ��,  ����@  �~(W���  ���   ����~ �|'/t��������R�P���  �Pd�����  �xd����(V���   ZY�t$�V���D�����[^_ÐUWVS��   ��  �Ʃ  ��@  ���   ��x;��  �  ���C(P�l$U���  �Pd�,$���  ���   �ǃ����  �|/t6��������R�T$U���  �Pl����t���T$R�W���  �Pd���{��tb�����   W���  ���   ����t7���  �pd��U���   ZYW�P�֋��   ����t	��U�Ѓ��    �Ĝ   [^_]Ív ���   ��x�;��  }����  �pd��U���   ��XY�?������   P�R�f�� �����$  ������������   P���������f��!�����������PU���  �Pd���{�������c����v UWVS��,�R  ��  �|$@�t$D��@  �E ���C  ���  ���[  �L$H��p������T$����L$�T$L���������1�T$��jh   @h,  h�  �LQ�L$ �TR�PT��jh����h,  h�  �t$,V�|$$W���  �RT��h����jh�  VW���  �R@��h����jh�  ��,  RW���  �R@��h����h,  jVW���  �R@��h����h,  jV���  R���  �R@�|$(��
��jh����jj�V
RW���  �RT�t$4���� h   ���6���RV�D$�PR���  �RDh   ��URV�D$$�P2R���  �RD��h�   hfff��U(RV�D$$���   R���  �RH�t$4��(�� �}��  �D$
   ��   ��j�P�D$h|  VW���  �R@��h����jh|  VW���  �R@��h����jh|  �D$�PW���  �R@�D$4��*�� 1���S����L$��E����L$�|$���g�v �L$�D$��jjW�D$�PRQj ������ h   ��D$������   P�GP�D$��#P���  �PD�D$�D$�����L$9�td�t$��   9��  ~R9��   u'��h�׳�jhz  �G�P�D$$��P���  �P@�� �6�0����$  ���C����L$�>���f��D$��  �}��   �L$�D$���   h   ���8���RW�t$�VR���  �RD�D$$�   �t$��<�$����jh�   P�D$ V���  �R@��h   �jh�   �D$PV���  �R@�� h   ����   RW�t$�VAR���  �RD���L$��jh����jj<Q�L$ �|$$���   R���  �RT�t$4��  �� h   ���>���RV��  R���  �RDXZjh�z �jj<�L$Q��@  R���  �RT���  �RD�� �}t<������j�PV�D$O  P�҃��   ��,[^_]�f��D$   ��   �G���f���������1���,[^_]�f��  ��k	  ��@  � ��t1����  ����Ív UWVS���  ��<	  �T$8��@  ���tg�D$0-�  ��9�S���  9�|I�|$4��,  ��;|$<7��,  ;t$<|+�p	9���   �p(9�|)�w	;t$<} �w;t$<|�����f��   ��[^_]Ív �q�t$N�
  ��   ��|  9�|�o(9l$<|v�;t$<|n�T$<)�����������   x�9��  ~�9��   ��   ���   �|$u�k�0��$   �x���PP���  ���   R���   R�Pd���V���f���  ���   9�},��6  9�|"9t$<�0�����  ;l$<|�    �������?  9��
���|  9������9t$<�������  ;|$<������������������   �����k�0��$   u�|$ �>����у����   P�4���������S���   ��W  ��@  ���t�|$tn�|$
t�{t�   ��[Ív ���e�����v �����  ���   R���   ���|$t0�L$�Q���^w���>��L$���   Ƅ�    �f��    뗅�~�Ƅ�    뉋$Ë$Ë$Ë<$Ë4$�  t���`������������������4����������T���t���`������������������4����������T���t���`������������������4����������T���New Open Save  * Length:  /home Open File Untitled.txt New.txt Save As TextEdit Quit [FW] cm_init: Done.
 fs_new_folder fs_new_file <Menu name=" </Menu> <Item label=" id=" <key> </key> <string> </string> CamelMenuDef [FW] Loading config for:  / Info.clist [FW] Picker Refresh...
 [FW] Picker Refresh Done.
 . [FW] Dialog Init...
 [FW] Dialog Init Done.
 ^ Name: Cancel    [FW] WARNING: cm_init called twice!
    [FW] cm_init: Setting up framework...
  [FW] Failed to allocate config buffer
  [FW] Config not found (or empty):   [FW] Config loaded successfully.
   %   2      #       *   &      )      $      	                %   /                        0   .         '   
                !                                         (          -                                                                          1      ,              "                                           +       %         	   �AZ �  ��
#  0@  pB�  �PU  B   �  �   @                     
                                                     !   "   &   '   (   )               *   +   ,   /   1       2�?���!wp���Lʽ|����h#���bϐ����+g=��!_^�tz5ӝ���rMw9J/q|aI�q���b*�|EI�%+R��	�P�Y�^47(2ӏigs2I��W>�i��*)��� c��Wm+�c%14t��hjі����"U+y��}Sn7���K��	9�xy��Bd8��iB����s!�Ql
7            TextEdit                                   �����  X          Untitled.txt                                                                                                                    �  �  �   �
  �H    �      O                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (,  ���o�-     �R     �O  
   �           �U     @               ���o                                                           �  �  �    �  �H  @    �  �  {     �  L  8     )     s    �  �&  %     B  �  [     0  �?   	    N     k       P  O     �   P  y        �   |     �   0  �     t  �  �     �   �(  �     �  �H       n  �  3    �   �  �     2   "  �    X  h  :     )  �  �     �   �
  �    �  D  |     �  `2       [  �  V     �  �  N     �   h  4     �   @	  D    \   x  d     S  D  �     ~  $       �  h   �    �  �  �     g   �  �       �  v     J  �  l    ;  �  D     �   �  t            �     
  �  \     (  T  �    2  �&  �    �  D  �     
    �    J  ,  :     j  T  5     �  `?          x  �     C   �  ~      on_file_picked_open on_file_picked_save on_paint cm_dialog_render doc_insert doc_backspace doc_delete get_visual_pos_of_index get_index_from_visual_pos ensure_visible move_vertical move_word on_input cm_dialog_input file_open_action cm_dialog_open file_save_action cm_dialog_save file_new_action on_mouse cm_dialog_click menu_cb cdl_main cm_init cm_dialog_init my_memcmp my_strstr my_strchr actions action_count config_count cm_bind_action execute_action_by_id internal_menu_callback strncpy_safe parse_menus_from_string parse_plist_xml cm_get_config cm_load_app_config cm_apply_menus cm_draw_image cm_draw_image_clipped cm_picker_refresh cm_picker cm_dialog_up_dir cm_dialog_select_dir cm_dialog_submit cm_dialog_handle_mouse  0     0     0     0     0     0     0     0     �       0�             T      �  2   �  j   E   1-  	S   X   r   r   r   r   r    2int z  
�   �   �   r    �  �   �   �   r   r   r    �  �   �   �   r   r    0�   d   �    �  #   
    2    
  3  
  )  2    4 	X  �   
X   �  4h  �  	r   � 
  h  2    
�   x  2        )  �		  �     �  4  �  M  c  ]  Y  c  �   w     !�  n  "�  �  %�     &�  $�  '�  (^  (�  ,8  )w  0Y  *�  4Q   +w  8w   .,  <   /P  @�  0o  D�  1�  Hi  2�  Lh  3�  Px  4�  T  5  X�  88  \�   9X  `q  :m  d   ;�  hs  <�  l�   =�  p�  >�  t  ?�  x*  @X  |�  A�  �J  B  �  C  �2  F$  ��  G$  �  H$  ��  IC  �J  J$  �    M�  ��   Na  �"  O  ��  P  ��  Q�  �<   R�  �h  S�  ��  T  �   U3  ��  VQ  �  W�  ��  X�  ��  [c  �        	  E   -  -   �    E   M  E   -   9  ]  E    R  5b  r   w     h  r   �       |  �  �  r      �  r   �    �  r    �  r   �    E   r    �  r   �    r    �  9   ,    r   r   G   y   �      P  r   r   r   r   r    1  o  r   r     r    U  �  r   r     r   r    t  �  r   r      �  �  r   r   r   r      �  �  r   r   r   r   r   r    �    9     r   �    x  �  8  E   r   -   #  R  E   R  -   W  6=  m  �     ]  �  �    -   r  r   �      -   �  �  �    r    �  �  �       �  r   �  �     �  -       �    r   �   
  7&     >  >  >  >   r   )  r   a  r   r   r    H  r     r   R  r    f  r   �  r   R  -  r   R  r    �  r   �  r   R  -  r    �  r   �  r   E   -  r   E   >   �  r     r   E   -  r      r   3  r    $  r   Q  �  �  �   8  ~  ]�  $_	�  �   _     _'E        _3b  ,`	�  �   `   +   `)r    �   `6r   $8  `R�  ( �  �   `]�  �  V  �     
  �  2    
  	  2   ? sys �  X2  �  �  T2  �   r   P2  �  �  �/  3   r   L2  �  r   H2  �  r   D2    r   t/  z  r   p/    r   �  !r   l/  Q  ��  @/  %J  �	   &*  �	  �     �r   
  r   r   r   r    '  ;8
          �   'Q  :W
        �   �   Gr   {
  r   r   r   r    (A   �r   �
  r    8�  ��  �  l  �  api �'�  V&*  �
  �   %J  �
   y  �
  ��}win �E   W;	  �  @0   
    2   � 
x  #  2    9  �F  )  r   )�  r    :�  m�  �   �P  *x r         *y r   $       btn m!r   �  �r   �  r   r   r   r    ;�  @   +  %  vr   6   4   �  wr   B   @   �  xr   R   L   �  {r   �   �   �  |r   �   �   *  F   �  �	  l  c  y  P  �  m   <�  kP  O   �=+  b>\  ah  4   ��  �  8
   �   Y�   |   ��  +[  Y  �  '  O    �   ��  +[  O  � len R	r   �   �    �    s  ��  x r   � y r   �w !r   �h (r   �bx 	r   �   �   by r   `  Z  2  
�  ��~%  	r   �  �  E  	r   �  �  cx 	r   �  �  cy r   $    �  	r   H  B  h  r   j  d  �	  ?	r   �  �  �   A
�  ��~num B
X  ��}�   Gr   7  r   r   r   r       �  i  r   �  �     c $  �  �  �  D   t 0%�  ��~   '   �  �  8r   @2  ,w  w  <  W
  ,m  u  
  �  2   � 
  �  2    ?  �B  @key �r   (A   �r     r    �  �	r   ;  �r   alt �r   A6  i �r    Bi �r     @  �@	  D  �n  dir �r   � �	  �   <  ��  t   ��  dir �r   � �  �	r   �hh  �r   �lC�  �	r   $  �	r   �  �  `  �	r       �    +	  F  6	  �    B  �P  y   �F  cx �	r   �hcy �r   �lE  �	r       v     D�  Yr   x  �   �  �   Y#r   � $  Y1r   �	cx Z	r   I  9  	cy [	r   �  �  <  \	r   �  �  [   ]	r   �  �  W   	i `r      �  �   �  _   dr   !     l   	c w  1  )     �  A�  �   ��  E�  A"r   h  `  �  A3>  �m  A?>  �	cx B	r   �  �  	cy C	r   �  �  2   	i Gr   �  �  B   	c H          �  5x  d   ��  �     	i 7r   Y  U     �  -  k   �	  /     	i /r   n  l    �  $�  ~   �E  c $  � �     	i &r   z  v    -�  �
  �  �e  !�  � "  "  "  F�  �
   �   �[  #�  �  �  �   $  �T$  �X$  �\.6  �   �  /7  �  �  F  n   .'  �   �  /,  #    f  n   s  �  �  �  �  	  y  �  �  n  �  n  �  B  �  B  -  	  B  	  N  	    �
  {
   -c  �  �   ��  Gc  �   �   bF  
   H#  �  [   �!1  � !;  �I#  �   �   ��  #1  O  M  #;  Z  X   �  c  �  P  �  m    �   �  4�  �      T    b  �  2   �  j   E   5-  	S   X   r   r   r   r   r    6int z  
�   �   �   r    �  �   �   �   r   r   r    �  �   �   �   r   r    0   d       �  #   
    2    
  7  
  ,  2     ]  �   
]   �  4m  �  	r   � 
  m  2    
�   }  2        ,  �	D  �  T   �  o  �  �  c  �  Y  �  �   �     !�  n  "�  �  %     &  $�  '!  (^  (:  ,8  )�  0Y  *�  4Q   +�  8w   .g  <   /�  @�  0�  D�  1�  Hi  2�  Lh  3  Px  45  T  5Y  X�  8s  \�   9�  `q  :�  d   ;�  hs  <�  l�   =�  p�  >�  t  ?  x*  @�  |�  A,  �J  B@  �  CU  �2  F_  ��  G_  �  H_  ��  I~  �J  J_  �    M  ��   N�  �"  O�  ��  P�  ��  Q�  �<   R
  �h  S7  ��  TZ  �   Un  ��  V�  �  W  ��  X  ��  [�  � O  O     D  E   h  h   �  Y  E   �  E   h   t  �  E    �  8�  r   �  O   �  r   �  O  O   �  �  �  r      �  r     O  �  r    �  r   !  O  E   r      r   :  O  r    &  9   g  O  r   r   G   y   �    ?  �  r   r   r   r   r    l  �  r   r   O  r    �  �  r   r   O  r   r    �  �  r   r   O   �    r   r   r   r   O   �  5  r   r   r   r   r   r      T  9   T  r   �    }  :  s  E   r   h   ^  �  E   �  h   �  9x  �  �  O   �  �  �  O  h   �  r   �  O  O  h   �  �  �  O  r    �  �    O  O   �  r   ,  �  O  :   h  @  O   1  U  r   �   E  ;&   Z  y  y  y  y   r   d  r   �  r   r   r    �  r   �  r   �  r    �  r   �  r   �  h  r   �  r    �  r   
  r   �  h  r    �  r   7  r   E   h  r   E   y     r   Z  r   E   h  r    <  r   n  r    _  r   �  �  �  �   s  ~  ]�  �  �   T  0-�  �   .�   

  /r   (�  0r   , 
  �  2   '  �	  2  	r    �
  	r   2  
  U  
�	  (A   
�	  ��
  !
�	  �W
  $	r   �9  %	r   �8  (�  �d	  1�	  �<a  2	r   � 
  �	  2    
  �	  2   ? 
  �	  2    
�  �	  2   ? 	  3�  =�	  6�	  �	  �  �  �	  
  �  �  &   >sys �   O  $2	I
  &id 3  �
  4�    A	  5)
  
I
  e
  2    }  7U
  �H  e
  8r   �H  
}  �
  2    6	  :�
   K  	  ;r   �J   >�
  &key ?  �  @
�
    
  �
  2   � ,
  A�
  
�
    2    �
  C�
  �?  H  Dr   `?  ?�	  O`2   A   �r   �(  �   ��  key �r   � �  }  len �r   s  o   )  �      fr   �&  �  ��  	  fr   � 	z  f$r   �mx f/r   �my f7r   �x i	r   �  �  y j	r     �  �	  u	r   C  ?  �	  v	r   n  h  fy �	r   �  �  s  }  idx zr   �  �  �  {r   �  �  ~(  �  �(  �   !�  �&  ]  i�  �  �  �   !�  '  h  j�  �       Z'  #   @�  Er   �&  %   �  mx E r   � my E(r   �btn E0r   �  �   �r   "  �  ��  	`  �r   � 	�
  �%r   �	  �0r   �	z  �;r   �x �	r       y �	r   z  r  �	  	r   �  �  �	  	r   �  �  
  	r   �  �  A�  	r   fy 0	r   	  	  "5$  �   S  i r   G	  ?	  R  idx r   k	  g	  iy  r   �	  z	  L
  (O  �	  �	  �$  ^    !�  I"  <  �v  �  �	  �	   '�  a"  G  ��  �	  �	    (�  �h   �  ��  ~  �
�	  ��~len �	r   �	  �	  �!  �   #�  ��  {   �#  	 	  �'O  � len �	r   
  
  B[   w `      C�	  �=  )len �r    D  ��  \   ��  2  �!O  
  
  �  �4O  /
  +
  	�  �KO  �	�
  �eO  �cb �~�  �  �   #Q  �0  �   �  	2  �!O  � 	�  �4O  �	�
  �KO  �cb �d�  ��     EJ  ��  V   �(�	  [�  3  ��  F@d�  y	  e�   �  f&   (�
  g&   ,�  h�	  0*uid i�	  1�  j�	  2*gid k�	  3
  l�  4 G  m4  	  o	r   D
  @
  �  p�  a
  W
  �  O  u	r   �
  �
    i wr   �
  �
    

  {r   �
  �
  �  �r       &  i  �  �r   +  '  �
  �r   =  ;   �  F   idx �r   G  E      
&   �  2    +�
  Hh  :   �^  "
  H&
  S  O  �   H8O  n  d  x HBr   �  �  y HIr   �  �  dw HPr   �dh HXr   �cx H`r   �cy Hhr   �cw Hpr   � ch Hxr   �$,�  -��  +f  E,  :   ��  �  E
  �  �  �   E2O  �  �  x E<r       y ECr   -  )  	�	  EJr   �	�	  EUr   �,c  -��  #r
  "�  D   �  	�
  "E   �  $�
  �r   T  �  �o  P  �$O  Ve  
�	  ��~)len r   �  
�  V�  	r   P $�	  �O  �  v   ��  key �'O  � �  O   i �r   A  =    %  ��  �  �2  xml �$�  � ptr ��  Y  Q  �   �	  ��  �  x  u  ��  �  �  �     w  �r   �  �  i �r   �  �  �  ��  	      ��      �     �
  ��  4  ,  �  �r   W  S  Q
  ��  r  f  �	  ��  �  �  "�  H   �  k �r   �  �   "d  L   �  k �r        �  �  :  �  W  �   �  �     �  .  �    %p  �  �  �j  buf ��      ptr ��  &  "    �  ��  7  5  :
  ��  C  ?  A  ��  T  R    �  �@'
  �r   `  \  m  ��  �  �  �
  ��  �  �  �
  ��  �  �  �
  �r   �  �  ~  �  �  �  �  �  �  j  �  �    �  "  �  �  j  �  �    Hl	  �L  8   ��  I�	  ��      src �+O  H  >  n �4r   y  o  i �	r   �  �   J*  m�  .�	  m!r   .t  m/r   Kid }O   /O	  cD  |   �2  id c'O  � �   i dr   �  �    %V  \�  N   �c  �  \!O  � �
  \3�  � /*  HD  �   ��  api H�  �  �  �  Ir   �J   0�  &�  $     ��  s &O  �  �  c &$r        $  �  �  �   �X  �	  O  � /	  3O  �Q  	r       �  	r   ,  (  �  8   i  r   ?  ;    X    0�  r   T  5   ��  s1 �  � s2 +�  �n =h  �p1 O  Q  O  p2 O  Z  X  Z  &   i h  i  a    L�  r   �  Mval !r    N�  �  �   �z  1�  � 1�  �2�  �  �  O�  4   4     mg  �  �  �  �  �  �  3�  C  �     �  +  �   P#  D  �   �31  '#  w   1  �1  21      �         I   :!;9I8   !I  H }  'I  '   :;9I  4 :!;9I  	4 :!;9I�B  
I  ! I/  4 :!;9I�B  4 :!;9I�B  4 :!;9I   :!;9I  U  4 :!;9I�B  :!;9  .?:!;9!'I<    .?:!;9!'@z   :!;9I  $ >     4 :!;9I  4 :!;9I  4 :!;9I  .?:!;9!'@|  U  4 :!;9I   :!;9I   .?:!;9!@z  ! 1  "4 1  # 1�B  $4 1  %.?:!;!�9!<  &.?:!;!�9!'<  '.?:!;9!'<  (.?:!;9!'I<  ) :!;!�9I  * :!;!�9I�B  + :!;9!&I  ,H }�  -.1@|  .1U  /4 1�B  0%  1   2$ >  3& I  4:;9  5 '  6&   7 'I  8.?:;9'I@|  9.?:;9'   :.?:;9'@z  ;  <. ?:;9@|  =. ?:;9   >.?:;9@z  ?.?:;9'   @ :;9I  A  B  C4 :;9I  D.?:;9'I@z  E :;9I�B  F1R�BUXYW  G 1R�BUXYW  H.1@  I1R�BUXYW    I   :;9I8   !I  H }  'I  '  4 :!;9I�B  4 :!;9I�B  	 :!;9I  
I  ! I/   :!;9I  4 :!;9I�B   :;9I  4 :!;9I�B  $ >  U   1�B   :!;9I�B   :!;9I8   :!;9I   :!;9I�B  U   :!;9I  :;9  4 :!;9I?  4 :!;9I  4 :!;9I     :!;9I�B  :;9!	   .?:!;9!'I@|  !1R�BUX!YW  "  #.?:!;9!'@|  $.?:!;9'I@|  %.?:!;9!'@|  & :!;9!
I8!   '1R�BUX!YW  (.?:!;9!@|  )4 :!;9!	I  * :!;9!I8  +.?:!;9!'@z  ,H}�  -I ~  . :!;9I  /.?:!;9!'@  0.?:!;9'I@z  1 1  24 1�B  34 1  4%  5   6$ >  7& I  8 '  9&   :   ; 'I  < :;9I8  =4 :;9I?<  >4 :;9I  ?4 G:;9  @.?:;9'I@z  A4 :;9I  BH }�  C.?:;9   D.?:;9'@  E. ?:;9@|  F:;9  G :;9I  H.?:;9'@z  I :;9I�B  J.?:;9'   K4 :;9I  L.:;9'I   M :;9I  N.1@z  O1R�BXYW  P.1@|   _            ��� ��W     �����V  ��(�  ��wv�      ��v D2  "(���Q��v D2  "(�  ��<�  ��v D2  "(<<#
�     JkPktP2                       ��P����}����}��� #P���P����}��� #P���� #����P����}��� #����
� #���
�� #��       ��W��
�#��
��#�         ��P����}��
��}�
���}         ��Q����}��
�@��
���}          ��:���W��:���W��:���W�
�:�       ��:r ���U�
�:r �      ��	����	��}�
�	��      ��	����	��}�
�	��         �	�	wh��	�	P�	�
wh��
�
wx�     ��0���V       ��P����}��P  ��	v <ut"���v <ut":+( �   ��P     ��r@���
p/  @�           ��:���Q��:���Q��Q��:���Q��:�        ��:���S��S��:�     ��R��R          ���� ���U��U��U���� �        ��0���P��P��0�   ��V        ��w p "��w p "��w p "1��w p "         ��� ��S��� ��S       ��:���R��:���R��R��:�        ��:���Q��Q��:�        ��0���P��P��0�          ��u p "��u p "1��u p "��u p "1��u p "     ��P��H2     ��U     ��P���h                    ��V��� ��V��� ��V��� ��V��� ��V��V       ��0���:v ���;v ���:v �       ��0���:v ���;v ���:v �  ��0�  ��3� �
            �/�/P�0�0P                   �+�,P�,�,
� 
�1&��,�,P�,�-
� 
�1&��-�.P�.�.p�}��.�.
� 
�1&��.�.P�.�.
� 
�1&�        �+�+
�
,1&��+�+w 1&��+�,
�
,1&��,�.
�
,1&�    �,�-�
,1&#(��.�.�
,1&#(�      �,�,ȟ�,�,V�.�.ȟ   �-�.V    �,�-	�u D��.�.	�u D�         �,�,
r P3  "��,�-R�-�-T3  �.�.R    �+�+� 
���+�+P �+�+�
,�             �"�"Q�"�#�H�#�%�D� "��%�*�
�1&� "��*�*�D� "��*�*�
�1&� "�         �"�"R�"�$�T�$�*�
,1&�"��*�*�
,1&�"�         �$�&V�&�*�T#(��*�*V�*�*�T#(�    �$�%ȟ�*�*ȟ    �%�*D��*�*D�         �'�(Q�(�)�L�)�*�T#���*�*�T#��        �%�&0��&�&�D�&�&P�&�(�D     �&�&V�&�(V            �&�&w~��&�&wj��'�'w~��'�'P�'�'���'�'w~�   �&�&Q �!�!�
�� �"�"�
,�         ��P��W�!�!P�!�!W   ��P     ��� ���      ������    ��@���@�         ��P��V���X���X��V             ��P��R���L���L��P��R          ��0����D��R���D��0�       ��w 1���W��W    ��0���0�     ��P���\   ��P   ��Q     ��� ���            �����S�����S���       �����R��R     �����Q     ��� ���            �����S�����S���       �����R��R     �����Q    ��0���S        ��S��S������S           ��U��P��U���\��U       ��P��V��V       ��S��	�J  1���S      ��0���P��0�     ��P���@     ��V�	�	V         ��	V�	�	v{��	�	P�	�V     ��	U�	�U          �	�	P�
�
P�
�
p��
�
q��
�
q p "#��
�q p "#�        �
�
P�
�
p��
�
q��
�
q p "#��
�
q p "#�    �
�
0��
�P    �
�
0��
�
P   ���     ��P��P   ��P     ��P��V   ��P  ��p v ���p v O-( �   ��P       ��V��P��V     ��P��R       ��p v ���r v ���u�v �-( ���r v �-( �           ��� ��Q��� ��Q���            �����V�����V���           �����S�����S���      ��0���P��P    ��0���U       ��� ��� ���      ��� ��P     �����Q     ozPz�W     ��P��U    ��0���V  5�   5�      0�p � �	p � #�*p � �      ��p 0r 8$"K  "���p 0� 8$"K  "����0� 8$"K  "�   ��R���  ��e�           ��P��p���P��P��P��R��P                  T                     T            �         ������ ���� ����	 ������ �������� �������� �������� ���� ���� ���� ���� ���� ���� �         ���� ������ ������ ��	�	� ���� ���� ���� ���� ���� �!�!�!�" �"�"�"�" �%�&�&�' �+�+�+�+ �+�+�+�+ �,�-�.�.�.�. �/�/�0�0 ^    @   �         L   U   h   	   	   x   �   ,     �!	f J fK�u	uf,	����"'�0�,g!	fK
 tug/�=  o+�<K	f���",	��.< <h .j ��t< <i $k ��t< <i &.K�	�	��?"g	f ��x+	��" � �K=[�# JK  �% 1 � f X �<( n   �d6 �* JL?�=  X( w   �f<J X- �	K$	�K,	�!��% f��' H� ' � � ��~<=	f  J � u �0 f> , X YYt�2K����	f# J f  K0 @ , X  Y�t2K��h�	f# J �  K*   < f4 tB 0 X  Yf$K��FP!	 $ Jg i�	*W�<0 v   J	K tK=	[0 v   JJ J g � gv�= Y.	uW;�	g	  �! g	d�N	+VWt	.K f]< c  	Mg: fgK/t=Z c   J#: a� �=   YJr�$�X�<iK"h�! �/ * <�<1 JP ? <: Jg J  ��Y1f	��!z<	Xi�vgY�1!e	�f# J- E �1 J f1 JE �h Xr E  r �1 .$ < � JF tP $  P �$ .��u	r� J'  v+ . f+ .@ t J � .A "p A Jf JA p �+ . J " x�JZ	 f�z�	���	f � f$ �"(  + ( �5 J �K JU (  U �( .d<�Y2H�$.f% XRJ/$& �" kf " f/ �G �" Q �" . �5 v% 
�! �  J � 5 z% �! �  J �( Xgt���q� �' �z< f% �/   � f+ �5 )�<��~% �6 ��� ��[�Y�	 fs	 �	ug	�, �9 :-u�!%�26�@D�LP�SPf{&ZZ" X$ �fqt$ f$ . </ J	uy<)��tw t	g�	m�<	Y<	Yf% �9 X# �6 X$ u8 X"t/	�	K	Y X	Y a	Y	rS   f> H . 	Y,A�	g �g tL)�#ZK ��1��YYY�/ t  �    <   �         �   �   �   �   x   �   @ T  g	 "     	Y.< J& * <1I/;h! ��K�g	  X.! �  	�f � �t& yX5'��	�	K
 s4!./��	h�����f�/I	r. J . J� qJJ@���Y<f&J�K .�g+h�	 t# f  	u u�" J" p X9�i]^ J�r;<X��	sf�<nf	
�D7k� ' �/ # <   J <+ J/=  	-.=  )7 ���x'��	!<P	��X	/	�	�u>!f�(�11<-h8) - 1I1. J1 X['<�<K��fN�-�<h�"/ ��Ju�!{Y�: $ : < � : t�CG : I$ : J* � �w< $ < < �K?C < I$ < J+ �< � �	J<P2�Y�!�tg�#%1�
�	[<S	�	�	�#	�  �1 	>!	�	�K	��.	�	�#	� �0 	?!	!	�<.�1J��y<z�2. i .�A<  ,;�!	 �# �  	�&tf �7 t> �Js/5��. �K �� f. tv� ��!�"/{L��f��	s�;  S �	�	fgx<.	l�<	f�'�!	f JKf	KL\Xgf J <  J J JK  = |=gf J <  J J JK  = <!�	f�@)��"L	 ���	t<	� �	�2	zd<0 J�= b  �Y,�/J.K+�)� cf J J !v��f�j���g�?Jf< � � � ff�f�<fgf�h���u� J�� t�� t��!uu z� � ���!K� t  f J �= ;KL!	 �s�- � <9 �   + . J
Z%Zu }+ .g J t	�&	Y &-.0<�� t9 t ��)� ��Y�L�' J�K �/ t J, <	u��	| Xu%� � yf/f% t�
f	s�f+ J�%� �h. �	m�8��M<t�t	g��<B��� � f��|��|�	 �.��|��|�	 �.x�M'����J�J$�&	u	I[����
 �E . � J	�w:�	�) pX J J <	�	�	���@X�	@2E� � �	�	���#��('*"� � f���0 O� .�+ ��� .5��� J�;OY�L�{��{�.��{� J fH�{�." �6 f, fi< � <( J" <: f0 <	gYF );XN�t	s[$  f	F( @G f8 .	gfX	[f .��*iS t4 <�.Vft��	if2 J f7 JO �C f	g	gjf1 � X6 �N �B f9 c� �0 s
�0<��E<tf'���LyyxfX	p�u	]<f	��t, XY-�-�	p	g. J: 
 ping close strncpy cdl_symbol_t menu_def_t version is_dirty send cm_dialog_input fs_exists min_diff label win_handle_t create_window cdl_exports_t stats doc_len target_x on_file_picked_save socket memcpy cm_dialog_render strncmp lib_name file_picker_cb_t symbol_count set_window_menu on_input ta_y memmove title fs_delete ensure_visible exports fs_rename free cur_y get_launch_args kernel_api_t sendto preferred_cur_x exec target_idx doc_backspace net_get_interface_info malloc memset mouse_cb_t ctrl fs_list process_events cm_dialog_save cm_dialog_click file_save_action move_vertical cm_dialog_init exit fs_create draw_image_scaled input_cb_t draw_text_clipped line_h sprintf cdl_main fs_read get_visual_pos_of_index print uint32_t item_count file_new_action menu_cb_t mem_total itoa win_w dns_resolve target_y paint_cb_t symbols move_word strlen cm_dialog_open new_idx recvfrom strcpy draw_rect_rounded item get_kbd_state blink doc_delete out_x realloc action_id on_mouse GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection snap_y doc_insert exec_with_args menu_cb func_ptr draw_rect cm_init get_ticks best_idx ta_h get_fs_generation file_open_action out_y strcmp win_h current_path doc_buffer http_get get_index_from_visual_pos mem_used draw_text scroll_y connect click_x click_y recv on_paint cursor_idx show_save_prompt fs_write bind on_file_picked_open shift key_content_end hlen cm_bind_action clist_path parse_plist_xml file_buf my_memcmp my_strchr cm_dialog_select_dir perm visible_items start_dir long long int cm_dialog_submit show long long unsigned int dates my_strstr parse_menus_from_string active selected_index config_count current_dir entry_count val_tag name_ptr full_path value attr initialized real_idx nlen default_name menu_end key_tag size short unsigned int i_idx cm_dialog_handle_mouse dirname max_read file_picker_t temp_menu_count needle temp_menus action_bind_t execute_action_by_id entries strncpy_safe filename id_p req_h haystack dest menu_idx cm_picker menu_tag req_w cm_dialog_up_dir cm_get_config list_h cm_picker_refresh list_y unsigned char is_dir item_h short int buff klen config_pair_t key_content_start icon lbl_p scroll_offset action_count cm_apply_menus func mode val_content_start vlen cm_load_app_config item_tag cm_draw_image_clipped win_handle flen win_y filter filter_ext val_content_end item_ptr key_name raw_entry_t internal_menu_callback filename_input app_bundle_path win_x cm_draw_image item_idx actions safe_div2 usr/apps/textedit_cdl.c /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/apps usr/apps/../../sys usr/apps/../lib cdl_defs.h camel_framework.h usr/lib/camel_framework.c usr/lib usr/lib/../../sys     ���� |�  L           �   A�A�AdEBA FEFA LWAG jAA�A� X       �   |   A�A�A\A FEFFA JAAG VA
A�A�DCBA L �        s  A�A�A�A�F�v�E�B�G�G�G�F�E�B�G�K�G�d�B�B�B�B�A�A�V�E�G�A�K�J�A�B�B�B�B�A�K�L�E�G�A�K�J�A�B�B�B�B�A�M�L�E�G�A�M�J�A�G�E�L�S�A�A�M�i�K�A�G�X���G�E�D�G�J�L���E�B�B�K�J�E�Z�E�B�G�S�G�F�E�F�M�A�G�E�J�A�A�E�N�A�D�D�L�G�G�G�G�H�F
A�A�A�A�CL�A�G�A�G�C�E�8       �  ~   A�A�A�A�AtA�A�A�A� 4         k   A�A�A�A�c�A�A�A�   (       x  d   A�A�A�^�A�A�4       �  �   A�A�A�A�y
�A�A�A�DP       x  �   A�A�A�A�C�
A�A�A�A�Dq
A�A�A�A�A<       P  y   A�A�A�C$P(E,F0\ xA�A�A�   $       �  t   A�BE��i�A�A� <       @	  D  A�A�A�A�C0�
A�A�A�A�C  �       �
  �  A�A�A�A�C<P@H0E4E8E<E@E0z
A�A�A�A�Bk<B@H0N<B@H0V<B@H0Z<B@H0J<B@H0P<B@H0P<B@H0R<A@H0K<B@T0(       h  4   A�CQGGG HA� t       �  �   A�A�CRG LGA LEFFA VA
A�A�CCBA LEF G$G(G,G0HAA�A�       P  O   C~G FH       �  �   A�A�A�jAAF HA
�A�A�DYgA ^   4       �  [   A�Cm
A�BH
A�CQ
A�B  �       �  l  A�A�A�F�]�L�E�E�B�A�L�C�A�K�A�E�E�Z�K�F�F�F�E�E�G�N�G�G�T�A�G�D�J�A�G�D�J�A�G�D�J�A�G�G�O�B�A�A�UA�A�A�C����C�A�G�       f)            j)            n)            r)        ���� |�  ,   �  T  5   A�A�k
�A�BC�A�   l   �  �  �   A�A�A�A�C0^<D@O<D@O0a4A8D<A@H0K
A�A�A�A�CGA�A�A�A�     �  $     D   �  D  �   A�ClG EEBF @A�B�W
A�DCA�0   �  �  N   A�A�AZJM VAA�A�X   �  D  |   A�A�A�A�C0|8D<A@L0W
A�A�A�A�ECA�A�A�A�T   �  �  �   A�Cl
A�CCW HC
A�BCG HC
A�BCG HCA�,   �  L  8   A�A�k
�A�BF�A�   �   �  �  �  A�A�A�A�CTaXB\K`NP}XD\A`NPKXD\A`JPgXK\A`LPAXD\A`NPiXG\A`JPGXK\A`JP�
A�A�A�A�A(   �    �  A�BF�����A�A�A�X   �  �  v   A�A�A�A�C0w8D<G@L0O
A�A�A�A�DEA�A�A�A��   �  T  �  A�A�A�A�F�Y�e�A�A�E�Z�N�G�C�K�L�A�G�A�G�C�W�I�E�B�A�L�E�A�A�L�K�A�e�K
A�A�A�A�BC�G�m�H
A�A�A�A�AC�M�E�,   �  �  D   A�ClAGA FCA�     �  ,  :   A�t
�CA�   �  h  :   A�t
�CA��   �  �  3  A�A�A�A�CLRPQ@_LEPH@IDEHBLAPLDBHALDPN@@HDLAPF@]HDLKPF@~HALTP[@bLAPo@C
A�A�A�A�DCLAP\@MHALJPL@  4   �  �  V   A�A�CX EKBG ]A�A� d   �  0  �   A�A�A�A�C z(A,D0N G(A,D0N G(A,G0]A�A�A�A�B ����  D   �  �  \   A�A�ASDDD U[
A�A�DAA�A�   X   �  D  �   A�A�A�A�C(R,J0L G,A0O m
A�A�A�A�AO(A,D0L  T   �  �  {   A�A�A�NJ ONGC LLD GADC JA�A�A�   �   �  h   �  A�A�A�A�F�j�D�E�]�R�G�E�L�G�E�C�L�J�G�O�P�A�G�A�A�C�K�G�A�E�L
A�A�A�A�D^
�A�I�A�P�C�DZ�H�J�M�G�A�L�     �  "  �  A�A�A�A�C@`HBLEPETEXE\I`FHBLEPETEXE\E`LLEPBTEXA\A`LLEPBTEXG\A`LLEPETBXA\A`LLEPETBXA\G`SHBLEPBTBXD\A`S@EDGHALHPNTDXA\H`LLEPETDXA\K`S@ZLBPATIXA\A`LLEPBTEXA\A`LLEPBTEXG\A`S@lHBLBPATHXA\B`H@EDQHDLHPW@eLEPBTEXD\H`L@JDGHALHPbTEXA\E`LLEPBTEXE\A`L@EDGHALHPL@GHBLEPBTBXA\O`V@EDGHALGPJLAHBLEPBTBXE\G`U@NDAHALJPE@H
A�A�A�A�CaA�A�A�A�   �  �&  %   T   �  �&  �  A�A�A�A�C0�
A�A�A�A�Dy4A8N<G@F0�<H@H0(   �  �(  �   A�Cs
A�DOM I    �  f)        �  j)        �  n)        �  v)        �  r)                                 ��   X2          T2          P2       '   �/  �     4   H2       ?   D2       H   L2       Q   t/       W   p/       ]   @2       e   l/       u   @0       }   @/  ,     �            �   �         �   �         �   �         �   �         �   �         �   �         �   �         �   $         �   T         �   4         �   t         �            ��    O       �   �J       �   �J       �    K                    ��  v)          r)        4  O       	 =  f)        S  j)        i  n)           0        �    �    �  �(  �     �  "  �    �  �H       �  �&  %     �  �  N     �  �  ~       L  8       P  y        `?       -  x  d     8  $       B  �  3    T  ,  :     b  h   �    s  �  \     �  �  [     �  D  �     �  �  �    �  �  �     �  �   |     �  0  �     �  �  t     �  P  O     �  �
  �    �  h  :       �  �     +  D  �     <  �  v     J  �  �     [  �&  �    k  �H  @    s  x  �     �  �  �     �  D  |     �  T  �    �  `2       �    s    �  �?   	    �  h  4     �  �  l    �  @	  D    �  �  V       �  D       �  {     )  T  5     3  �  �     J    k     X      �      textedit_cdl.c sys doc_buffer doc_len current_path cursor_idx scroll_y is_dirty win_w win_h blink.1 preferred_cur_x menus.0 exports .L183 .L201 .L203 .L193 .L192 .L191 .L190 .L189 .L188 .L187 .L186 .L184 camel_framework.c initialized.0 temp_menu_count temp_menus __x86.get_pc_thunk.si __x86.get_pc_thunk.di _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.dx __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ parse_plist_xml cm_dialog_input cm_dialog_render action_count cm_dialog_handle_mouse cm_bind_action doc_insert strncpy_safe ensure_visible config_count doc_delete my_strchr cm_picker_refresh cm_draw_image cm_dialog_submit cm_dialog_save menu_cb cm_init parse_menus_from_string on_mouse on_file_picked_save cm_dialog_open move_vertical file_new_action on_input cm_draw_image_clipped get_visual_pos_of_index cm_dialog_up_dir cm_get_config file_save_action cm_dialog_click actions get_index_from_visual_pos my_strstr execute_action_by_id cm_load_app_config cm_picker on_paint file_open_action cdl_main move_word cm_dialog_init cm_apply_menus cm_dialog_select_dir my_memcmp internal_menu_callback doc_backspace on_file_picked_open  .symtab .strtab .shstrtab .text .rodata .gnu.hash .data .got .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_rnglists .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                          z)                 !         |)  |9  �                 -         (,  (<  d  
             )   ���o   �-  �=  �  
             3         @/  @?  �                   9          0   @                    >          0   @                   G         @0  ,@  �                  L         O  _  �                U         �O  �_                 ]         �R  �b  �                 e              �e  �-                 q              ��  �	                               T�  D                 �              ��  @                  �              خ  �                 �              f�  �                 �      0       _�  �                �      0       ��  �                 �              ��  X                 �   	      �U  �e  @   
                           �  �     (         	              ��  l                               �  �                  