ELF              D   4   x(      4    (                 �  �                    �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �D$D$Ív �D$+D$Ív �D$�D$�f��L$��t�D$����1�Ð�D$�Ѓ��f�S���.   ���  �D$��t� ��t����k���R�Ѓ��������[Ë$�Math Library Initialized!
                                                        ��q         ���`�T}G�T��TV��17�T                        CamelMath                             `                      add                                 sub                                mul                                div                             $   is_even                         8                        �   ���o�           �  
   ;            T     0               ���o                                                           2   D   7     
      	           
        $        %   8   
            	      math_add math_sub math_mul math_div math_is_even cdl_main  H     �     �     �     �          &
       �             {       �  1   =  �   C   �   	P   U   o   o   o   o   o    int �  
�   �   �   o    u  �   �   �   o   o   o    �  �   �   �   o   o    
0�     �    �  #       	1    A      #  	1     	R  �  
R   (  4b    	o   �   b  	1    �   r  	1    �   #  
�	  �     &  -  �  F  v  V  �  \  �   p  �  !�  �  "�  �  %�   =  &�  $N  '�  (�   (�  ,T   )p  0�  *�  4Y  +p  8.  .%  <�  /I  @8   0h  D�  1�  H�  2�  L  3�  P�   4�  T(   5  X�  81  \�  9Q  `&  :f  d�  ;�  hi  <�  l  =�  pM   >�  t}   ?�  x   @Q  |F  A�  �  B�  �  C  ��  F  �P  G  �V  H  ��  I<  �k   J  �!  M�  ��  NZ  �	  Ox  �-  Px  ��   Q�  �<  R�  �{  S�  �p  T  �J  U,  �    VJ  ��   W�  ��   X�  �  [\  �          C   &  &   8    C   F  C   &   2  V  C    K  [  o   p     a  o   �       u  �  �  o      �  o   �    �  o    �  o   �    C   o    �  o   �    o    �  8   %    o   o   E   v   �    �  I  o   o   o   o   o    *  h  o   o     o    N  �  o   o     o   o    m  �  o   o      �  �  o   o   o   o      �  �  o   o   o   o   o   o    �    8     o   �    r  �  1  C   o   &     K  C   K  &   P  6  f  �     V  �  �    &   k  o   �      &   �  �  �    o    �  �  �       �  o   �  �     �  &  �     �    o   �     &     7  7  7  7   o   "  o   Z  o   o   o    A  o   x  o   K  o    _  o   �  o   K  &  o   K  o    }  o   �  o   K  &  o    �  o   �  o   C   &  o   C   7   �  o     o   C   &  o    �  o   ,  o      o   J  �  �  �   1  �   ]}  
$_	{  �  _   �   _'C     c  _3Z  
,`	�  �  `   5  `)o    �   `6o   $0  `R�  ( {    `]�  �  O  p  �  {  �  	1    -  %�  `  B   -�        6�  D   7   �@	  api 6'�  �  ^   o   8   
   �g	  num o   �  `  o   $      ��	  a o   � b o   � �  o      
   ��	  a o   � b o   � �  o      	   ��	  a o   � b o   � �  o       	   �a o   � b o   �   I   :!;9I8   !I  'I  '   :!;9I   :!;9I  I  	! I/  
:!;9  .?:!;9!'I@z  $ >  4 :!;9I  %     $ >  & I  :;9   '  &       'I  4 :;9I  .?:;9'I@|  .?:;9'I@z                    {           �     7   �         C   K         ]        
�L�L�>KM�11 �,</ J .	K� g net_get_interface_info memmove cdl_main set_window_menu draw_text my_exports strchr fs_delete math_is_even get_fs_generation strstr http_get draw_rect_rounded fs_create win_handle_t kernel_api_t symbol_count sendto func_ptr paint_cb_t menu_def_t dns_resolve strlen bind itoa cdl_exports_t ping strcpy my_symbols long unsigned int close mem_used fs_exists cdl_symbol_t recv mouse_cb_t strncpy get_kbd_state math_mul memset exec_with_args draw_image get_ticks realloc input_cb_t draw_text_clipped exec action_id get_launch_args item_count process_events items create_window send char sprintf fs_list mem_total math_div strcmp k_api free recvfrom draw_rect menu_cb_t print GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection memcpy exit math_add socket uint32_t fs_rename math_sub lib_name fs_read label strncmp draw_image_scaled malloc connect version fs_write usr/lib/math.c /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/lib usr/lib/../../sys cdl_defs.h      ���� |�             	             	             
          $             8   
   $       D   7   A�C\G EIA�       {                                  ��      ,        `  �                  ��            '   {         =           S      
     \   $        e   8   
     r       	     {   D   7     �      	      math.c my_exports my_symbols _DYNAMIC __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ math_mul math_div math_is_even math_add cdl_main math_sub  .symtab .strtab .shstrtab .text .rodata .gnu.hash .data .got.plt .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_aranges .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                                             !      2                         -         �   �  0                )   ���o   �   �  <                3               �                   9                              B               �   	             K         �  �  p   	            S             ;                  [              �  *
                 g              �  T                 u                                   �              "  �                  �      0       �  F                �      0       B%  h                 �              �%  �                  �   	      T  T  0                              H&  �               	              ('  �                                �'  �                  