ELF              �  4   ,.      4    (                 d  d           ,  ,  ,  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      S���  �ÿ  ��`   ��t,���   ���T$���`   ���   =�� w�D$�    ��[�f����L$���[�f�S���J  ��c  ��X�������	)Ѝ�����	)��Љ������)Ѝ��90  ��X������   1���Ӌ�`   ���   �d   1����w���C��[�f�WVS��   ���  ��`   ����   ��8   ��   ��u&���V(�v �    �@   ��9�u�ǃ      ��   �+�������   @�
   �����   ��8   �V(1���9�u����  �gfff�������)�[^_�f��d   [^_Ív 1�[^_�f��   3  �T$��`   ��x���Ë$Ë$Ë$�                                               a          xR�����l����                 90                              SysMon                                �                      cpu                             �   ram                                 ,                                                                                                            �  ���o�          �  
   G            L                    ���o                                                              \   v     >   �       )   �   �            Z      sysmon_get_ram_usage calculate_cpu_load sysmon_get_cpu_usage cdl_main  h     �     �     �
       �             �      �  1   �  H   C   "  	P   U   o   o   o   o   o    int �  
�   �   �   o    E  �   �   �   o   o   o    �  �   �   �   o   o    
0�   B   �    v  #       1    -      #  1     	R  �   
R   �  4b  �  	o   �   b  1    �   r  1        #  
�	  �     7  -  n  F  �   V  g  \     p  �  !�  �   "�  �  %�   �  &�  $P  '�  (l  (�  ,�   )p  0�   *�  48   +p  8`   .%  <�  /I  @<  0h  D�  1�  H�  2�  Lv  3�  PN  4�  T�   5  X>  81  \�   9Q  `G  :f  d   ;�  h  <�  l�   =�  p�  >�  t,  ?�  x�   @Q  |�  A�  �7  B�  �  C  ��  F  �3  G  �  H  �`  I<  ��  J  �    M�  ��   NZ  ��  Ox  �F  Px  �  Q�  �3   R�  �>  S�  �N  T  �   U,  �   VJ  �  W�  �#  X�  �X  [\  �          C   &  &   �    C   F  C   &   2  V  C    K  [  o   p     a  o   �       u  �  �  o      �  o   �    �  o    �  o   �    C   o    �  o   �    o    �  8   %    o   o   E   v   �    �  I  o   o   o   o   o    *  h  o   o     o    N  �  o   o     o   o    m  �  o   o      �  �  o   o   o   o      �  �  o   o   o   o   o   o    �    8     o   �    r  �  1  C   o   &     K  C   K  &   P  6  f  �     V  �  �    &   k  o   �      &   �  �  �    o    �  �  �       �  o   �  �     �  &  �     �    o   �     &     7  7  7  7   o   "  o   Z  o   o   o    A  o   x  o   K  o    _  o   �  o   K  &  o   K  o    }  o   �  o   K  &  o    �  o   �  o   C   &  o   C   7   �  o     o   C   &  o    �  o   ,  o      o   J  �  �  �   1    ]}  
$_	{  �   _   �  _'C        _3Z  
,`	�  �   `   +   `)o    �   `6o   $   `R�  ( {  n   `]�  �  O  sys �  (  o   �  1   	 	  �     	m  	o   �  	x  
o   �  {  >	  1    	|   9.	  �  	�  >�  @  �  B�  �     ��	  api B'�  �  S  2    Z   ��	  �  %�	  � �  8�	  � &   �  o   
  sum *	o   avg -	o   �	  i !o     i +o     !�   o   \   v   �_
  	2  1      "h  	o   �  o         U   o   .   *    #�	  �   �   ��	  D   B   �	  $�	       �
  �	   %�	  I     �
  &   �	  S   M   �	  n   j   '�	     �	  �   �      (1  
     I   :!;9I8   !I  'I  '   :!;9I  I  ! I/  	4 :!;9I  
:!;9  4 :!;9I  4 1�B  $ >   :!;!29I  4 :!;9!	I�B  4 1  %     $ >  & I  :;9   '  &       'I  4 :;9I  .?:;9'I@z   :;9I  .?:;9'@|  .?:;9I        !.?:;9I@|  "4 :;9I  #.1@z  $1  %1R�BUXYW  &U  '1U  (H }   �               ��R��S��p{�     ��p d���R  ��0�      ��0���Q��Q    ��q :���q :�  ��0�                  �                   ���� ���� �    7   �         E   M         _   B     1�	fK' f�fg t# �) r�Wt�'
ti&<	Xifg' � X  >=J>��f+ !: ' f + : ' t 	u�f X=#t�i	r 	�' /+ # . v	��1 d X nt.,f�	� g ping close strncpy cdl_symbol_t menu_def_t version send fs_exists label win_handle_t tick_delta create_window cdl_exports_t my_symbols calculate_cpu_load socket memcpy strncmp lib_name symbol_count set_window_menu memmove fs_delete fs_rename free get_launch_args kernel_api_t sendto exec net_get_interface_info malloc memset mouse_cb_t fs_list process_events exit fs_create draw_image_scaled draw_image input_cb_t draw_text_clipped my_exports sprintf strchr cdl_main fs_read used_mb print uint32_t item_count menu_cb_t mem_total itoa dns_resolve paint_cb_t char seed strlen recvfrom strcpy draw_rect_rounded get_kbd_state realloc action_id spike GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection exec_with_args sysmon_get_cpu_usage func_ptr long unsigned int draw_rect get_ticks items get_fs_generation cpu_samples strcmp http_get strstr mem_used draw_text connect recv sysmon_get_ram_usage base sample_idx initialized fs_write total_mb bind usr/lib/sysmon.c /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/lib usr/lib/../../sys cdl_defs.h     ���� |�  (           Z   A�CD
A�CLA�         \   v   A�CpA�H       �   �   A�A�A��
�A�A�CF
�A�A�DC�A�A�         �            �            �            �                                 ��
   (                        (     !   �       -   �       8   @  ,     C   �  H                  ��N   �        d   ,        m   �        �   �        �   �        �   �   �     �   \   v     �       Z     �   �        sysmon.c sys seed.0 cpu_samples initialized sample_idx my_exports my_symbols __x86.get_pc_thunk.cx _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ sysmon_get_cpu_usage calculate_cpu_load sysmon_get_ram_usage cdl_main  .symtab .strtab .shstrtab .text .gnu.hash .data .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_rnglists .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                          �                 %         �  �  (                !   ���o   �  �  0                +               �                   1         �  �                   :         �  �  L                   ?         ,  ,  �   	             H         �  �  P   	            P             G                  X              d  �
                 d              S                   r              m!  �                  �              �!                     �              "  "                  �              ?"  �                 �      0       6$  �                �      0       �)  j                 �              <*  �                  �   	      L  L                                (+  0              	              X,  �                                M-  �                  