ELF                 4   \�      4    (                  R   R           \  L  L  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      UWVS��(�  ��P%  �|$@h��t$L�t$LW�t$L���	  �P@���   �D$(� ���   �G�D$,�Ǎ��  �� �D$0���D$�; th����SW�t$���	  �RD����Q��
9�uڋD$� �   �����	D�����	  h � �j
j���   � ����L$$�P���   ��	���L$L�DP�R@�� ��[^_]Ív UWVS���  ��h$  ���   �D$�Í��  �݃�QRjPSU���	  �R`�EP ��9�u�PjPj �D$�  P���	  �P\���   �    ��,[^_]�f�UWVS���F  �#  �D$�t$0���ta���   ���   ���   �D$�"����OI�Y������\$؈���t'F�E ��
u�@�E �    ��~�\$�������uك�[^_]�@�E �    ��	�   1�뢈T$�\$������E ��Y�T$뇐S���  ��?#  ��d���P�)���X������������p����$������[�f�WVS�Z  ��#  �D$D$uD���   ���  PjPj S���	  �P\��Q��9�u獆�   �     ���   �     ���h���[^_�UWVS����  �Ơ"  ������U������_X��s���P��D   W���	  �Pl�����  ����x���PW���	  �Pl����ty����~���PW���	  �Pl�����  ��������PW���	  �Pl������   ��W���	  ���   ����ta��������P������<$������,$��������=���   ���  QjPj S���	  �P\��Q��9�u獆�   �     ���   �     ���H�����$   �     P���	  h�   j W�P\����[^_]Ív �������P�Q�����빃�������P�=���Z�������1����������$�#�����X����$�������z�������	  �@��[^_]��f�WVS�F  ���   �D$��
��   ��tP�P���^wD��$   ���~7�r�1��D   ����   ���O���   �6�z�9����������[^_Í�$   ���~�H���D   � ���   ���~�J����   � ���������� �f�����[^_Ív WVS��   �  ��.   ��$  ���	  ���   ���  �����	  RjPj S�P\��Q��9�u��h   �\$S���	  �PY_������P��d���W���	  �Pd�$���	  ���   �܅���   ��SW���	  �Pd�������$�������<$�����������$�s��������%�����j ������������h,  h�  ������P���	  �P<�Ã�������P���  W���	  �PdXZ������P�GP���	  �Pdǆ�	     ������jWS���	  �PX��$�����   [^_Ív ��������P����������S���f��VS�t$��t&�D$�T$��f�@B9�t��8�t���)�[^Ð1�[^Ív UWVS����  �À  �t$0��tr�L$4��tj���t$<���&  ���   ��Z�t$@���&  ���   ��)�x=1��ŉ|$��v F�D$9�'�|$0�PU�t$<W�Q�������uމ����[^_]�f�1���[^_]ËD$�L$��u	�f�9�t
@���u�1�ÐS���  ���  �D$���"  ��uoǃ�"     ���&  ��������R���h@  j ���������&  �P\��$   �     ��  �     ǃ�"      ���&  �������T$ � ��[����t� ��t�������T$��[��f���[Ív VSR�j    ��$   ���0�����&  �t$�ҍ�D   ��P�Qd����L$$�L� @���X[^�f�UWVS���  ���  �D$0�D$��$   ���~N��D   �D$��1��
f�E��$9.~4���t$W���&  �Pl����u��D� �T$�D� ��t��[^_]���v ��[^_]�S���  ��O  �T$�D$��dt@��etS��x9��"  ��[�f������ ����D���"  P�1�������[Ð�������P��������[Ð�������P��������[ÐVS�L$�t$�\$1����f��@9�t���u��� [^Ð�� [^�UWVS��@��  �  �D$�\$Tǀ�"      h   j ���"  �|$(W�ǋ��&  �P\���; �5  ���� ����|$$��&����D$(��"  �D$�f��]�} �  ���t$,S�\$�z����Ń�����  ���t$0P���^�������t��p���"  ����  �S���"  �P����  �����D$�1��f�F@�T����t
��"t��u����߉\$ ؋L$� ���\$��-���PU������D$ �����M  9��4�����5����D$߉l$,�f��D$��8�   ���D$9��  ���t$ V�\$�����ƃ�����   9D$��   �D$��8�   ����   ����;���PV�R���������um���\$��C���PV�5����������p����P���e����D- �(���D$ ËD$�1���v ���?���@�T�T���.�����"u��$����P��t��\- ����D$ ËD$�1��@�T�T���b�����"�Y�����u��O����l$,�]�} �������<[^_]�1��n���U��WVS��L�H  ���  �E��  �M��    �8 ��  ��H����}���f����M���$  �}���E�� �B	�z	 �b  ���u�P���������K  ���u�P����������4  �p����N���PV����������  W��)��~�   �E�RV�}�W�q���Y^��U���R�E�P����������   ���u�P����������   �p����^���PV�j���������   �Eċ ���(����U���W�����M��P���&  �Pd���U���)�=�   ~��   �U�PV�Eċ �����M��D P�����XZ��h���PW���&  �Pl�����U���������Eċ �����M��D P�������U�������e�[^_]�UWVS���  ��0  ��  ���~N1�1ۍ�$  �D$�f�C��   9~1���t$8�D$�P���&  �Pl����u׋D$�D ��[^_]Ív 1���[^_]�f�UWVS��   �  �õ  ��$�   ��u���P���&  ��4$���&  ��������,$���&  �_XV�|$W���&  �Pd�<$���&  ���   ����~�|�/t��������R�P���&  �Pd�����&  �pd��W���   ZY������R�P���$   ���&  �P�ƃ�����   Ph   j V���&  �P\��h�  VW���&  �P ����~>� ��V�����4$���&  �P���&  ��(����$����   �Č   [^_]Ð�������P���&  ��<$���&  ��,$���&  ����&  �4$�P��1��Č   [^_]Ã����&  ������R���1��܍v S���u  '  �L$���&  ��t#��t���"  ��~������S���"  PQ�RX����[�S�4  �  �\$�T$�L$���&  ��t�@L��t�\$�L$�T$[���[�f�S��  �  �\$�T$�L$���&  ��t�@L��t�\$�L$�T$[���[�f�UWVS��8�  ��h  ������P���&  ����&  ������  ��
  �|$Ǉ�      ��h   �P�ƃ����g  Ph   j V���&  �P\��j@V�G(P���&  �P(������  �D$    ���&  �������|$�������|$�t$�T$f��> ��   ���t$V�Pl������   �~0�����&  ��u7���t$�L$���   U�Pl�����  ���&  �L$���    ��   �L$���  ��?F�i�T$���  ��V�,	����T$���   Q�Pd�T$Չ�$  �F(��(  �����&  �D$�T$��@9T$�.����t$��V�P�D$ǀ�   ����ǀ�       ���&  �������$�����,[^_]Ív ��V���   �D$,�,$���&  ���   ��9D$�y�����U�L$()��P���&  �Pl�����W������&  ���������&  �_����VS���  ��6  ���&  ������R������&  h   j ��
  V�P\�    ���&  �������$���[^�f�UWVS���2  ���  �D$ �l$$�|$(��
  �   �C    ���&  �Rd��tb��P�CP�ҋ��&  �@d����tX��U�S(R�Ћ��&  �@d����t6��W���   R�ЋD$<���   ƃ�    ���������[^_]Ð�� ���떍������������VSQ�z
  ��(  �t$�t$ �t$ �t$�t$�!�����
  �@   ����t���&  �t$�   �D$�BdZ[^��f�X[^�UWVS���&
  ���  ������S��
  �n(U���&  �Pl����t=��U���&  ���   ����~-�P��|'/u�E�Ht)�T(��/u��D( ���������[^_]�u�V)�����u���S�F(P���&  �Pd����f��D' ��1�븐WVS�v	  ��$  ����
  �~(W���&  ���   ����~ �|'/t��������R�P���&  �Pd�����&  �xd����(V���   ZY�t$�V���D�����[^_ÐUWVS��   ��  �ơ  ��
  ���   ��x;��  �  ���C(P�l$U���&  �Pd�,$���&  ���   �ǃ����  �|/t6��������R�T$U���&  �Pl����t���T$R�W���&  �Pd���{��tb�����   W���&  ���   ����t7���&  �pd��U���   ZYW�P�֋��   ����t	��U�Ѓ��    �Ĝ   [^_]Ív ���   ��x�;��  }����&  �pd��U���   ��XY�?������   P�R�f�� �����$  ������������   P���������f��!�����������PU���&  �Pd���{�������c����v UWVS��,�N  ���  �|$@�t$D��
  �E ���C  ���&  ���[  �L$H��p������T$����L$�T$L���������1�T$��jh   @h,  h�  �LQ�L$ �TR�PT��jh����h,  h�  �t$,V�|$$W���&  �RT��h����jh�  VW���&  �R@��h����jh�  ��,  RW���&  �R@��h����h,  jVW���&  �R@��h����h,  jV���  R���&  �R@�|$(��
��jh����jj�V
RW���&  �RT�t$4���� h   ���
���RV�D$�PR���&  �RDh   ��URV�D$$�P2R���&  �RD��h�   hfff��U(RV�D$$���   R���&  �RH�t$4��(�� �}��  �D$
   ��   ��j�P�D$h|  VW���&  �R@��h����jh|  VW���&  �R@��h����jh|  �D$�PW���&  �R@�D$4��*�� 1�������L$������L$�|$���g�v �L$�D$��jjW�D$�PRQj ������ h   ��D$������   P�GP�D$��#P���&  �PD�D$�D$�����L$9�td�t$��   9��  ~R9��   u'��h�׳�jhz  �G�P�D$$��P���&  �P@�� �6�0����$  ���C����L$�>���f��D$��  �}��   �L$�D$���   h   ������RW�t$�VR���&  �RD�D$$�   �t$��<�$����jh�   P�D$ V���&  �R@��h   �jh�   �D$PV���&  �R@�� h   ����   RW�t$�VAR���&  �RD���L$��jh����jj<Q�L$ �|$$���   R���&  �RT�t$4��  �� h   ������RV��  R���&  �RDXZjh�z �jj<�L$Q��@  R���&  �RT���&  �RD�� �}t<�� ���j�PV�D$O  P�҃��   ��,[^_]�f��D$   ��   �G���f��������1���,[^_]�f��  ��c	  ��
  � ��t1����&  ����Ív UWVS���  ��4	  �T$8��
  ���tg�D$0-�  ��9�S���  9�|I�|$4��,  ��;|$<7��,  ;t$<|+�p	9���   �p(9�|)�w	;t$<} �w;t$<|�����f��   ��[^_]Ív �q�t$N�
  ��   ��|  9�|�o(9l$<|v�;t$<|n�T$<)�����������   x�9��  ~�9��   ��   ���   �|$u�k�0��$   �x���PP���&  ���   R���   R�Pd���V���f���  ���   9�},��6  9�|"9t$<�0�����  ;l$<|�    �������?  9��
���|  9������9t$<�������  ;|$<������������������   �����k�0��$   u�|$ �>����у����   P�4���������S���   ��O  ��
  ���t�|$tn�|$
t�{t�   ��[Ív ���e�����v �����&  ���   R���   ���|$t0�L$�Q���^w���>��L$���   Ƅ�    �f��    뗅�~�Ƅ�    뉋$Ë$Ë4$Ë$Ë<$�  user@camel: $  help clear exit ls Listing  :
  Command not found:  /home Directory changed to:  Camel OS Terminal v1.0
 Terminal Shell Clear [FW] cm_init: Done.
 fs_new_folder fs_new_file <Menu name=" </Menu> <Item label=" id=" <key> </key> <string> </string> CamelMenuDef [FW] Loading config for:  / Info.clist [FW] Picker Refresh...
 [FW] Picker Refresh Done.
 . * [FW] Dialog Init...
 [FW] Dialog Init Done.
 Open Save ^ Name: Cancel     Camel OS Terminal
 Commands: help, clear, ls, cd, exit
     (Directory listing not fully linked in this demo)
 [FW] WARNING: cm_init called twice!
    [FW] cm_init: Setting up framework...
  [FW] Failed to allocate config buffer
  [FW] Config not found (or empty):   [FW] Config loaded successfully.
   %   /             (         '      !          #             "   .             &           )   ,            +   $         	             
                                  %                                                                              *                            -                                    %             5Z�A� -&hC @ sL+�
H                        
                                                           #       %   '               (   )   *   -           2�?���Ƣ��!wp���Lʽ|����h#���bϐ x�tz5ӝ���rMw9J/q|aI�b*�|�b��EI�%�	�P�Y�^47(2ӎigs�u���(���+�f c��Wm+�c%1*��hjі����"�Cy���Rn7ө�1���K��	9�xy��Bd8��iB���YIE��    Terminal                        
                               /                                                                                                                               �$  @&  P  `  �E      	  L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �!  ���o #     |O     �L  
   i           �Q     8               ���o                                                           %  �	  �    �   �E  @    "   (&       �  0  {       �	  8            �     2  �  %     b   P  `     c  �<   	    r   �%  �     �  t  �     �   �  �     Y    �     �   �E       �  �  3    !  T  �    *   $&       �  �  :     �   `  �     �   �  |     �  `/       �    V     �   8  N     I     :        @&  �    �   �  �     2   �   n     �   h         �  �      	  �     {   �%       M     v     �      u    n  ,  D     
    &       j   �  �    �  ,  \     >   X  �     [  �  �    I    �    �  �  �     =  X  �    }  p  :     �   �  5     U   �$  �     �   `<        on_paint blink_state term_buffer cur_row cur_col term_scroll term_print term_prompt current_path menu_cb execute cmd_line cmd_pos on_input cdl_main my_memcmp my_strstr my_strchr cm_init actions action_count config_count cm_bind_action execute_action_by_id internal_menu_callback strncpy_safe parse_menus_from_string parse_plist_xml cm_get_config cm_load_app_config cm_apply_menus cm_draw_image cm_draw_image_clipped cm_picker_refresh cm_picker cm_dialog_init cm_dialog_open cm_dialog_save cm_dialog_up_dir cm_dialog_select_dir cm_dialog_submit cm_dialog_render cm_dialog_handle_mouse cm_dialog_click cm_dialog_input    @%     D%     H%     L%     P%     T%     X%     �       �  4           �      �  1   %  Q   C   /  	P   U   o   o   o   o   o    int �  
�   �   �   o    J  �   �   �   o   o   o    �  �   �   �   o   o    0�   K   �    �  #   	    1    y    	  #  1     	R  �   
R   �  4b  �  	o   � 	  b  1    	�   r  1        #  �	  )     <  -  y  F  �   V  �  \     p  �  !�  �   "�  �  %�   >  &�  $U  '�  (�  (�  ,�   )p  0�   *�  4A   +p  8^   .%  <�  /I  @  0h  D�  1�  H	
  2�  L�  3�  PY  4�  T�   5  XC  81  \�   9Q  `R  :f  d   ;�  h�  <�  l�   =�  p�  >�  t;  ?�  x�   @Q  |�  A�  �B  B�  �  C  ��  F  �  G  �	  H  �k  I<  ��  J  �    M�  �z   NZ  �G  Ox  �   Px  �  Q�  �3   R�  �I  S�  �0  T  �   U,  �%  VJ  �  W�  �  X�  �]  [\  �          C   &  &        C   F  C   &   2  V  C    K  [  o   p     a  o   �       u  �  �  o      �  o   �    �  o    �  o   �    C   o    �  o   �    o    �  8   %    o   o   E   v   �    �  I  o   o   o   o   o    *  h  o   o     o    N  �  o   o     o   o    m  �  o   o      �  �  o   o   o   o      �  �  o   o   o   o   o   o    �    8     o   �    r  �  1  C   o   &     K  C   K  &   P  6  f  �     V  �  �    &   k  o   �      &   �  �  �    o    �  �  �       �  o   �  �     �  &  �     �    o   �     &     7  7  7  7   o   "  o   Z  o   o   o    A  o   x  o   K  o    _  o   �  o   K  &  o   K  o    }  o   �  o   K  &  o    �  o   �  o   C   &  o   C   7   �  o     o   C   &  o    �  o   ,  o      o   J  �  �  �   1  �   ]}  $_	{  �   _   �  _'C        _3Z  ,`	�  �   `   +   `)o    �   `6o   $:  `R�  ( {  l   `]�  �  O  	  �  1     sys �  @/  	  	  1   1   P 
l  �  @&  
x  o   (&  
�  o   $&  
�  o    &  
8   �  �%  
  o   �%  
�  �  �$  �   ��  �$  !�  ��     u  �=
  api �'�  � �   �
=
  ��}win �C         �  �M
  @.  "   
  i �o   !       �  �  �  �  �  �  �  �  �  �   	  M
  1   � 	r  ]
  1     �  ��
  m �o   i �o   #i �o     $5  s    �   ��
  x so   � y so   �w s!o   �h s(o   �=   I   r xo   ,   *     �   [�
  key [o    %(  6�  �  ��  &�     (  i >o    �  �  s  �  {  �  �  �  �  �    �    �  '  �  5  �  C  �   '  0  :   ��  /  �  ;  �  I  �   ($   X  �   �	  )str    9   3   *   c "  X   P   �  	    	    +L  �   n   �;  �   0   y o   x   v     ,]
  P  `   ��  g
  � p
  �-]
  t  8   �g
  p
  .y
  t     �  /z
   �  �    0�
  `  �   ��
  �   �   1�
  �   �  D   [�  �
  �   �      �
    �   �  4�  s       �    �  �  2   %  Q   E   5/  	S   X   r   r   r   r   r    6int �  
�   �   �   r    J  �   �   �   r   r   r    �  �   �   �   r   r    0   K       �  #   
    2    y  7  
  ,  2     ]  �   
]   �  4m  �  	r   � 
  m  2    
�   }  2        ,  �	D  )  T   <  o  y  �  �   �  �  �     �  �  !�  �   "�  �  %   >  &  $U  '!  (�  (:  ,�   )�  0�   *�  4A   +�  8^   .g  <�  /�  @  0�  D�  1�  H	
  2�  L�  3  PY  45  T�   5Y  XC  8s  \�   9�  `R  :�  d   ;�  h�  <�  l�   =�  p�  >�  t;  ?  x�   @�  |�  A,  �B  B@  �  CU  ��  F_  �  G_  �	  H_  �k  I~  ��  J_  �    M  �z   N�  �G  O�  �   P�  �  Q�  �3   R
  �I  S7  �0  TZ  �   Un  �%  V�  �  W  �  X  �]  [�  � O  O     D  E   h  h      Y  E   �  E   h   t  �  E    �  8�  r   �  O   �  r   �  O  O   �  �  �  r      �  r     O  �  r    �  r   !  O  E   r      r   :  O  r    &  9   g  O  r   r   G   y   �    ?  �  r   r   r   r   r    l  �  r   r   O  r    �  �  r   r   O  r   r    �  �  r   r   O   �    r   r   r   r   O   �  5  r   r   r   r   r   r      T  9   T  r   �    }  :  s  E   r   h   ^  �  E   �  h   �  9x  �  �  O   �  �  �  O  h   �  r   �  O  O  h   �  �  �  O  r    �  �    O  O   �  r   ,  �  O  :   h  @  O   1  U  r   �   E  ;&   Z  y  y  y  y   r   d  r   �  r   r   r    �  r   �  r   �  r    �  r   �  r   �  h  r   �  r    �  r   
  r   �  h  r    �  r   7  r   E   h  r   E   y     r   Z  r   E   h  r    <  r   n  r    _  r   �  �  �  �   s  �   ]�  �  �  T  0-�  �   .�   ~  /r   (  0r   , 
  �  2   '  �	  Z  	r    	  	r   �  
  �  
�	  (�	   
�	  ��	  !
�	  ��  $	r   �q  %	r   ��	  (�  ��  1�	  �<�  2	r   � 
  �	  2    
  �	  2   ? 
  �	  2    
�  �	  2   ? X  3�  =  6�	  p      r  �  �  �  &   >sys �   L  $2	I
  &id 3  	  4�    �  5)
  
I
  e
  2    
  7U
  �E  �  8r   �E  
}  �
  2    �  :�
   H  n  ;r   �G   >�
  &key ?  �  @
�
    
  �
  2   � �  A�
  
�
    2    >	  C�
  �<  �  Dr   `<  ?�	  O`/   a  �r     �   ��  key �r   � �   }  len �r   �   �    G  �    �  fr     �  ��  	~	  fr   � 	s	  f$r   �mx f/r   �my f7r   �x i	r   �   �   y j	r   ]  U  i  u	r   �  �  P  v	r   �  �  fy �	r   �  �  �   }  idx zr   �  �  �  {r       �  �  �  �   !�  >  �   i�  �  E  A   !�  I  �   j�  �  ]  [   �  #   @0  Er   �  %   �  mx E r   � my E(r   �btn E0r   �  �  �r   T  �  ��  	 
  �r   � 	�	  �%r   �	~	  �0r   �	s	  �;r   �x �	r   x  l  y �	r   �  �  i  	r       P  	r   ?  ;  �  	r   V  R  A�  	r   fy 0	r   o  g  "y  �   S  i r   �  �  �   idx r   �  �  iy  r   �  �  �  (O      �  ^    !�  �  �   �v  �  !     '�  �  �   ��  2  0    (  ��  �  ��  �  �
�	  ��~len �	r   I  A    �   #�  �0  {   �#  	G  �'O  � len �	r   h  f  B�  w �     C1  �=  )len �r    D�  �,  \   ��  �  �!O  t  p  �  �4O  �  �  	�  �KO  �	�	  �eO  �cb �~�  �S  �   #~  �t  �   �  	�  �!O  � 	�  �4O  �	�	  �KO  �cb �d�  �     E�  �  V   �(W  [�  3  ��  F@d�  �  e�     f&   (+	  g&   ,�  h�	  0*uid i�	  1�  j�	  2*gid k�	  32  l�  4 G�	  m4  O  o	r   �  �  q  p�  �  �  �  �  u	r   �  �  t   i wr   $       ~  {r   R  L    �r   p  l  �   i  �  �r   �  �  y	  �r   �  �     F   idx �r   �  �      
&   �  2    +R	  H�  :   �^  �  H&
  �  �  �   H8O  �  �  x HBr   �  �  y HIr       dw HPr   �dh HXr   �cx H`r   �cy Hhr   �cw Hpr   � ch Hxr   �$,�  -��  +
  Ep  :   ��  q  E
  $     �   E2O  ?  5  x E<r   l  f  y ECr   �  �  	+  EJr   �	�  EUr   �,�  -��  #	  ",  D   �  	h	  "E   �  $6	  �r   �  �  �o  �	  �$O  V|  
�	  ��~)len r   �  
�  V  	r   P $B  �O     v   ��  key �'O  � 2  O   i �r   �  �    %B  ��	  �  �2  xml �$�  � ptr ��  �  �  >   "  ��  �  �  �  ��      N     
  �r   #    i �r   G  A    ��  c  _  �	  ��  w  s  ^     I	  ��  �  �  *  �r   �  �  �  ��  �  �  �  ��    	  "�  H   �  k �r   M  I   "�  L   �  k �r   a  ]   C  �  ~  �  �  �   �
  �   V
  �  r
  �    %�  �X  �  �j  buf ��  s  q  ptr ��  �  |  i   
  ��  �  �  �  ��  �  �  X  ��  �  �  �	  �  �@�  �r   �  �  �  ��  �  �  	  ��  �  �  �	  ��  	  	  1	  �r   	  	  �  �  �  �  �  �    j  1  �  H  �  f  �  �  j    �    H�  ��	  8   ��  I
  ��  q	  g	  src �+O  �	  �	  n �4r   �	  �	  i �	r    
  �	   J�	  m�  .  m!r   .
  m/r   Kid }O   /�  c�  |   �2  id c'O  � 3   i dr   
  
    %m  \8  N   �c  �  \!O  � 	  \3�  � /f  H�  �   ��  api H�  1
  +
  �  Ir   �G   0�  &�  h     ��  s &O  N
  J
  c &$r   b
  ^
   $8  �  �  �   �X    O  � �  3O  �h  	r   v
  r
  �  	r   �
  �
    8   i  r   �
  �
  G  X    0�  r   �  5   ��  s1 �  � s2 +�  �n =h  �p1 O  �
  �
  p2 O  �
  �
  �  &   i h  �
  �
    L%
  r   �  Mval !r    N�  	  �   �z  1�  � 1�  �2�  �
  �
  O�  x	   x	     mg  �  @  <  �  R  P  3�  �	  �   W	  �  o	  �   P#  �  �   �31  '#  �   �   ��   21  j  \  �         I   :!;9I8   !I  H }  'I  '   :!;9I  ! I/  	I  
4 :!;9I?   :!;9I  4 :!;9I�B  :!;9  $ >  4 :!;9I   :!;9I  .?:!;9!' !  4 :!;9!I     1   1   1�B  %     $ >  & I  :;9   '  &       'I   4 :;9I  !.?:;9'I@|  "U  #  $.?:;9'@|  %.?:;9@  &  '.?:;9@z  (.?:;9'@z  ) :;9I�B  *U  +.?:;9@|  ,.1@|  -1XYW  .1  /4 1  0.1@z  11R�BXYW    I   :;9I8   !I  H }  'I  '  4 :!;9I�B  4 :!;9I�B  	 :!;9I  
I  ! I/   :!;9I  4 :!;9I�B   :;9I  4 :!;9I�B  $ >  U   1�B   :!;9I�B   :!;9I8   :!;9I   :!;9I�B  U   :!;9I  :;9  4 :!;9I?  4 :!;9I  4 :!;9I     :!;9I�B  :;9!	   .?:!;9!'I@|  !1R�BUX!YW  "  #.?:!;9!'@|  $.?:!;9'I@|  %.?:!;9!'@|  & :!;9!
I8!   '1R�BUX!YW  (.?:!;9!@|  )4 :!;9!	I  * :!;9!I8  +.?:!;9!'@z  ,H}�  -I ~  . :!;9I  /.?:!;9!'@  0.?:!;9'I@z  1 1  24 1�B  34 1  4%  5   6$ >  7& I  8 '  9&   :   ; 'I  < :;9I8  =4 :;9I?<  >4 :;9I  ?4 G:;9  @.?:;9'I@z  A4 :;9I  BH }�  C.?:;9   D.?:;9'@  E. ?:;9@|  F:;9  G :;9I  H.?:;9'@z  I :;9I�B  J.?:;9'   K4 :;9I  L.:;9'I   M :;9I  N.1@z  O1R�BXYW  P.1@|   �             ��P��S  �
�
0�  =`0�     ��� ��V��V         ��R��R��R���_  ��0�           ��	� �	�	P�	�
� �
�
P�
�
�    �	�	�  �
            �/�/P�0�0P                   �+�,P�,�,
� 
�1&��,�,P�,�-
� 
�1&��-�.P�.�.p�}��.�.
� 
�1&��.�.P�.�.
� 
�1&�        �+�+
�
,1&��+�+w 1&��+�,
�
,1&��,�.
�
,1&�    �,�-�
,1&#(��.�.�
,1&#(�      �,�,ȟ�,�,V�.�.ȟ   �-�.V    �,�-	�u D��.�.	�u D�         �,�,
r P0  "��,�-R�-�-T0  �.�.R    �+�+� 
���+�+P �+�+�
,�             �"�"Q�"�#�H�#�%�D� "��%�*�
�1&� "��*�*�D� "��*�*�
�1&� "�         �"�"R�"�$�T�$�*�
,1&�"��*�*�
,1&�"�         �$�&V�&�*�T#(��*�*V�*�*�T#(�    �$�%ȟ�*�*ȟ    �%�*D��*�*D�         �'�(Q�(�)�L�)�*�T#���*�*�T#��        �%�&0��&�&�D�&�&P�&�(�D     �&�&V�&�(V            �&�&w~��&�&wj��'�'w~��'�'P�'�'���'�'w~�   �&�&Q �!�!�
�� �"�"�
,�         ��P��W�!�!P�!�!W   ��P     ��� ���      ������    ��@���@�         ��P��V���X���X��V             ��P��R���L���L��P��R          ��0����D��R���D��0�       ��w 1���W��W    ��0���0�     ��P���\   ��P   ��Q     ��� ���            �����S�����S���       �����R��R     �����Q     ��� ���            �����S�����S���       �����R��R     �����Q    ��0���S        ��S��S������S           ��U��P��U���\��U       ��P��V��V       ��S��	�G  1���S      ��0���P��0�     ��P���@     ��V�	�	V         ��	V�	�	v{��	�	P�	�V     ��	U�	�U          �	�	P�
�
P�
�
p��
�
q��
�
q p "#��
�q p "#�        �
�
P�
�
p��
�
q��
�
q p "#��
�
q p "#�    �
�
0��
�P    �
�
0��
�
P   ���     ��P��P   ��P     ��P��V   ��P  ��p v ���p v O-( �   ��P       ��V��P��V     ��P��R       ��p v ���r v ���u�v �-( ���r v �-( �           ��� ��Q��� ��Q���            �����V�����V���           �����S�����S���      ��0���P��P    ��0���U       ��� ��� ���      ��� ��P     �����Q     ozPz�W     ��P��U    ��0���V  5�   5�      0�p � �	p � #�*p � �      ��p 0r 8$"H  "���p 0� 8$"H  "����0� 8$"H  "�   ��R���  ��e�           ��P��p���P��P��P��R��P                  �              �       �            #         ������ �
�
�
�
 �         ���� ������ ������ ��	�	� ���� ���� ���� ���� ���� �!�!�!�" �"�"�"�" �%�&�&�' �+�+�+�+ �+�+�+�+ �,�-�.�.�.�. �/�/�0�0 �    7   �          L   U   =   =   h   +     � Y��	 v	�Y  d ��	Y<	f>�	�&t	����!	 	!0#( G yu�"��-
 �.)\<)-.�v	g	!;YJ g' X �fXz<J$g+  !�)<�廻�� t�( Z$ � 	��	�v�J!�	 �
� <
	t <
� <
� �	u�( k�$ � 	��	�u� f�	b�<! �; �	�yf	f<	ntJ!
�
X<qX1 & �	YX	��Y!)�-X�	oJ�K=��K=/	w�X,t�	g	  �$ b  � �[� �	���v-�Y�0�	rf �    <   �          �   �   {   {   h   �   @ �  g	 "     	Y.< J& * <1I/;h! ��K�g	  X.! �  	�f � �t& yX5'��	�	K
 s4!./��	h�����f�/I	r. J . J� qJJ@���Y<f&J�K .�g+h�	 t# f  	u u�" J" p X9�i]^ J�r;<X��	sf�<nf	
�D7k� ' �/ # <   J <+ J/=  	-.=  )7 ���x'��	!<P	��X	/	�	�u>!f�(�11<-h8) - 1I1. J1 X['<�<K��fN�-�<h�"/ ��Ju�!{Y�: $ : < � : t�CG : I$ : J* � �w< $ < < �K?C < I$ < J+ �< � �	J<P2�Y�!�tg�#%1�
�	[<S	�	�	�#	�  �1 	>!	�	�K	��.	�	�#	� �0 	?!	!	�<.�1J��y<z�2. i .�A<  ,;�!	 �# �  	�&tf �7 t> �Js/5��. �K �� f. tv� ��!�"/{L��f��	s�;  S �	�	fgx<.	l�<	f�'�!	f JKf	KL\Xgf J <  J J JK  = |=gf J <  J J JK  = <!�	f�@)��"L	 ���	t<	� �	�2	zd<0 J�= b  �Y,�/J.K+�)� cf J J !v��f�j���g�?Jf< � � � ff�f�<fgf�h���u� J�� t�� t��!uu z� � ���!K� t  f J �= ;KL!	 �s�- � <9 �   + . J
Z%Zu }+ .g J t	�&	Y &-.0<�� t9 t ��)� ��Y�L�' J�K �/ t J, <	u��	| Xu%� � yf/f% t�
f	s�f+ J�%� �h. �	m�8��M<t�t	g��<B��� � f��|��|�	 �.��|��|�	 �.x�M'����J�J$�&	u	I[����
 �E . � J	�w:�	�) pX J J <	�	�	���@X�	@2E� � �	�	���#��('*"� � f���0 O� .�+ ��� .5��� J�;OY�L�{��{�.��{� J fH�{�." �6 f, fi< � <( J" <: f0 <	gYF );XN�t	s[$  f	F( @G f8 .	gfX	[f .��*iS t4 <�.Vft��	if2 J f7 JO �C f	g	gjf1 � X6 �N �B f9 c� �0 s
�0<��E<tf'���LyyxfX	p�u	]<f	��t, XY-�-�	p	g. J: 
 ping close strncpy cdl_symbol_t menu_def_t version send cmd_line fs_exists label win_handle_t create_window cdl_exports_t socket memcpy strncmp lib_name symbol_count set_window_menu on_input memmove fs_delete exports fs_rename free get_launch_args kernel_api_t sendto cmd_pos exec term_prompt net_get_interface_info malloc memset mouse_cb_t fs_list process_events term_buffer cur_row exit fs_create draw_image_scaled input_cb_t draw_text_clipped sprintf cdl_main fs_read uint32_t item_count cur_col blink_state menu_cb_t mem_total itoa dns_resolve term_print paint_cb_t symbols strlen recvfrom strcpy draw_rect_rounded get_kbd_state realloc action_id GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection exec_with_args menu_cb func_ptr draw_rect get_ticks get_fs_generation strcmp current_path http_get mem_used draw_text connect execute recv on_paint fs_write bind term_scroll key_content_end hlen cm_bind_action clist_path parse_plist_xml file_buf my_memcmp my_strchr cm_dialog_select_dir file_picker_cb_t perm visible_items start_dir long long int cm_dialog_submit show long long unsigned int dates my_strstr parse_menus_from_string active cm_dialog_input selected_index config_count current_dir cm_dialog_save entry_count val_tag name_ptr full_path value attr initialized real_idx nlen default_name menu_end key_tag size short unsigned int i_idx cm_dialog_handle_mouse dirname max_read file_picker_t cm_init temp_menu_count cm_dialog_open needle temp_menus action_bind_t execute_action_by_id entries strncpy_safe cm_dialog_click filename title id_p req_h haystack dest menu_idx cm_picker menu_tag req_w cm_dialog_up_dir cm_get_config list_h cm_picker_refresh list_y unsigned char is_dir item_h short int buff klen config_pair_t key_content_start icon lbl_p scroll_offset action_count cm_dialog_render cm_dialog_init cm_apply_menus func mode val_content_start vlen cm_load_app_config item_tag cm_draw_image_clipped win_handle win_h flen win_w win_y filter filter_ext val_content_end item_ptr key_name raw_entry_t internal_menu_callback filename_input app_bundle_path win_x cm_draw_image item_idx actions safe_div2 /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/apps/terminal_cdl.c usr/apps usr/apps/../../sys cdl_defs.h usr/lib/camel_framework.c usr/lib usr/lib/../../sys camel_framework.h      ���� |�  l           �   A�A�A�A�C<T@DDDHALDPm0U4A8A<D@L0`<K@BDBHTLXPF0CA�A�A�A�T       �   n   A�A�A�A�C0c4B8A<A@P0E4B8B<J@XA�A�A�A�   <       X  �   A�A�A�A�C0|
A�A�A�A�A  $         :   A�CR FF VA�8       P  `   A�A�A�bBBA Od�A�A�  �       �  �  A�A�A�A�C,R0H,A(G,G0L K(G,A0L G(G,A0L K(G,A0L K,A0O G,G0X O$B(B,A0O p$K(B,A0F C
A�A�A�A�DC,G0H E,G0F,F0d RA�A�A�A�  8       `  �   A�A�A�j
�A�A�AJ�A�A��          u  A�A�A�F�n�B�B�A�I�G�E�E�J�A�G�G�Z�K�A�A�r�J�B�F�F�E�E�G�N�G�G�J�A�G�D�Y�B�A�A�UA�A�A�D����C�G�J�       �            �            �        ���� |�  ,   �  �  5   A�A�k
�A�BC�A�   l   �  �  �   A�A�A�A�C0^<D@O<D@O0a4A8D<A@H0K
A�A�A�A�CGA�A�A�A�     �  h     D   �  �  �   A�ClG EEBF @A�B�W
A�DCA�0   �  8  N   A�A�AZJM VAA�A�X   �  �  |   A�A�A�A�C0|8D<A@L0W
A�A�A�A�ECA�A�A�A�T   �  	  �   A�Cl
A�CCW HC
A�BCG HC
A�BCG HCA�,   �  �	  8   A�A�k
�A�BF�A�   �   �  �	  �  A�A�A�A�CTaXB\K`NP}XD\A`NPKXD\A`JPgXK\A`LPAXD\A`NPiXG\A`JPGXK\A`JP�
A�A�A�A�A(   �  X  �  A�BF�����A�A�A�X   �     v   A�A�A�A�C0w8D<G@L0O
A�A�A�A�DEA�A�A�A��   �  �  �  A�A�A�A�F�Y�e�A�A�E�Z�N�G�C�K�L�A�G�A�G�C�W�I�E�B�A�L�E�A�A�L�K�A�e�K
A�A�A�A�BC�G�m�H
A�A�A�A�AC�M�E�,   �  ,  D   A�ClAGA FCA�     �  p  :   A�t
�CA�   �  �  :   A�t
�CA��   �  �  3  A�A�A�A�CLRPQ@_LEPH@IDEHBLAPLDBHALDPN@@HDLAPF@]HDLKPF@~HALTP[@bLAPo@C
A�A�A�A�DCLAP\@MHALJPL@  4   �    V   A�A�CX EKBG ]A�A� d   �  t  �   A�A�A�A�C z(A,D0N G(A,D0N G(A,G0]A�A�A�A�B ����  D   �  ,  \   A�A�ASDDD U[
A�A�DAA�A�   X   �  �  �   A�A�A�A�C(R,J0L G,A0O m
A�A�A�A�AO(A,D0L  T   �  0  {   A�A�A�NJ ONGC LLD GADC JA�A�A�   �   �  �  �  A�A�A�A�F�j�D�E�]�R�G�E�L�G�E�C�L�J�G�O�P�A�G�A�A�C�K�G�A�E�L
A�A�A�A�D^
�A�I�A�P�C�DZ�H�J�M�G�A�L�     �  T  �  A�A�A�A�C@`HBLEPETEXE\I`FHBLEPETEXE\E`LLEPBTEXA\A`LLEPBTEXG\A`LLEPETBXA\A`LLEPETBXA\G`SHBLEPBTBXD\A`S@EDGHALHPNTDXA\H`LLEPETDXA\K`S@ZLBPATIXA\A`LLEPBTEXA\A`LLEPBTEXG\A`S@lHBLBPATHXA\B`H@EDQHDLHPW@eLEPBTEXD\H`L@JDGHALHPbTEXA\E`LLEPBTEXE\A`L@EDGHALHPL@GHBLEPBTBXA\O`V@EDGHALGPJLAHBLEPBTBXE\G`U@NDAHALJPE@H
A�A�A�A�CaA�A�A�A�   �  �  %   T   �    �  A�A�A�A�C0�
A�A�A�A�Dy4A8N<G@F0�<H@H0(   �    �   A�Cs
A�DOM I    �  �        �  �        �  �        �  �        �  �                                 ��   @/          @.          �$  ,     $            ��    L       6   �G       D   �G       T    H                    ��_   �        u   �        �   L       	 �   �        �   �        �   �        �   \%        �   X  �    �     �       �$  �       T  �    *  �E       7  �  %     N  8  N     ]  @&  �    i  �%       q  �	  8     ~  `<       �  h       �  �  3    �  p  :     �  �  �    �  ,  \     �  P  `     �  �%  �     �   &       �  �  �     �  �	  �        :       $&       &  t  �     5  `  �     >  �  :     T  X  �     _  �  �     p     v     ~    �    �  �E  @    �  �  �     �  �  |     �  �  �    �  `/       �  �  �    �      �     �  �<   	    �  (&       �     u    �  �   n          V       ,  D       0  {     3  �  5     =  	  �      terminal_cdl.c sys menus.0 exports camel_framework.c initialized.0 temp_menu_count temp_menus __x86.get_pc_thunk.si __x86.get_pc_thunk.di _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.dx __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ parse_plist_xml cm_dialog_input current_path cm_dialog_render action_count cm_dialog_handle_mouse cm_bind_action term_buffer cmd_pos strncpy_safe config_count my_strchr cm_picker_refresh cm_draw_image cm_dialog_submit cm_dialog_save menu_cb cmd_line blink_state cm_init parse_menus_from_string term_prompt cur_col cm_dialog_open on_input cm_draw_image_clipped term_print cm_dialog_up_dir cm_get_config cm_dialog_click actions my_strstr execute_action_by_id cm_load_app_config cm_picker execute on_paint cur_row cdl_main term_scroll cm_dialog_init cm_apply_menus cm_dialog_select_dir my_memcmp internal_menu_callback  .symtab .strtab .shstrtab .text .rodata .gnu.hash .data .got .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_rnglists .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                          �                 !      2   �  �.  �                -         �!  �1  X  
             )   ���o    #   3  |  
             3         �$  �4  �                   9         @%  @5                   >         \%  \5                   G         �%  h5  �&                  L         L  \  �                U         �L  �\  �              ]         |O  |_  i                 e               b  �&                 q              ƈ  �                               ��  �                 �              [�  @                  �              ��  �                  �              ��  u                 �      0       �  /
                �      0       1�  �                 �              �  0                 �   	      �Q  �a  8   
                           �                 	              �  T                               p�  �                  