ELF              \  4   �,      4    (                 �  �           x  x  x  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      UWVS���s  ��\  �l$0�|$4�\$8�L$<�L$�D$@�D$�T$D��   ����   ����   �T$��h   @QS�OQ�MQ�P@��   �� ��z ��T$�T$��Q�t$SWU�P@��h���@jSWU��   �P@���t$��   ���   �@�)É�������\$�������������T$��t@A��   �D$<�����|$�|$8�L$4�D$0�BD��[^_]���v ��V ��]���f���[^_]�U��WVS��,�M  ��:  �u�}�E�E��M�M�U�U܋U�U؋�   ����   ��h����Q�u�WV�P@����   �EԋU�R�u�M܅���   ��d��   �E��ȸ��Q�������)�PWV�M��Q@��h����j�u�WV��   �P@��h����j�u��M�D�PV��   �P@��h�����u�jWV��   �P@�� ��   �E�����M�M�E   �}�U��T��U�@@�e�[^_]���v �d   �N���f�1��E�����e�[^_]��     �T$��   ��x���Ë$Ë$Ë4$�                                            ��         ���M�5�V0p            CamelGUI                                                     btn                                 prog                               x                        �  ���o�     @        
   ,            l                    ���o                                                           #   \             <                 gui_draw_button gui_draw_progress cdl_main      @     d     �
       �             w      �  1   �  H   C   .  	P   U   o   o   o   o   o    int �  
�   �   �   o    D  �   �   �   o   o   o    	  �   �   �   o   o    
0�   B   �    �  #       	1    9      #  	1     	R  �   
R   �  4b  �  	o   �   b  	1    �   r  	1        #  
�	  �     6  -  }  F  �   V  {  \     p  �  !�  �   "�  �  %�   K  &�  $O  '�  (�  (�  ,�   )p  0�   *�  48   +p  8[   .%  <�  /I  @4  0h  D�  1�  H�  2�  L�  3�  PU  4�  T�   5  X=  81  \�   9Q  `N  :f  d   ;�  h  <�  l�   =�  p�  >�  t$  ?�  x�   @Q  |�  A�  �>  B�  �  C  ��  F  �+  G  �  H  �g  I<  ��  J  �    M�  ��   NZ  �T  Ox  �>  Px  �  Q�  �3   R�  �E  S�  �F  T  �   U,  �  VJ  �"  W�  �  X�  �W  [\  �          C   &  &   �    C   F  C   &   2  V  C    K  [  o   p     a  o   �       u  �  �  o      �  o   �    �  o    �  o   �    C   o    �  o   �    o    �  8   %    o   o   E   v   �    �  I  o   o   o   o   o    *  h  o   o     o    N  �  o   o     o   o    m  �  o   o      �  �  o   o   o   o      �  �  o   o   o   o   o   o    �    8     o   �    r  �  1  C   o   &     K  C   K  &   P  6  f  �     V  �  �    &   k  o   �      &   �  �  �    o    �  �  �       �  o   �  �     �  &  �     �    o   �     &     7  7  7  7   o   "  o   Z  o   o   o    A  o   x  o   K  o    _  o   �  o   K  &  o   K  o    }  o   �  o   K  &  o    �  o   �  o   C   &  o   C   7   �  o     o   C   &  o    �  o   ,  o      o   J  �  �  �   1    ]}  
$_	{  �   _   �  _'C        _3Z  
,`	�  �   `   +   `)o    �   `6o   $z   `R�  ( {  i   `]�  �  O  sys �  t  {  �  	1    w   9�     �  >�  �  �  B�  \     �G	  api B'�  �  �   )   <  ��	  x )o         y )#o   %   !   w )*o   :   6   h )1o   O   K     )8o   f   `   u  )J&   ��   0	o   �   �    f         �x o   �   �   y !o   �   �   w (o   �   �   h /o   �   �   B   >  ��  Io   �U   &       v   	o       tx !o   .  *  ty "o   @  >     I   :!;9I8   !I  'I  '   :!;9I   :!;9I�B  I  	! I/  
:!;9  $ >   :!;9I  4 :!;9I�B  4 :!;9I  4 :!;9!	I�B  %     $ >  & I  :;9   '  &       'I  4 :;9I  .?:;9'I@z   :;9I  .?:;9'@   :;9I�B  .?:;9'@   D            ��� ���      ������     ������     ������     ������T0+( d-( ����  �� �T0+( d-( �Xd�      �� ���       �����      �����      �����   Ls���x�   ��p 6�     ��P���    ��Q                  w          \    7   �         B   J         \   R     2	f�(�	P J�[/#  </.	�/t	�0 �    "f��JJ=sX�S�2	f�<�r�	��u�u<f�t<�=szX��,��	� g ping close strncpy cdl_symbol_t menu_def_t version send fs_exists label win_handle_t color create_window cdl_exports_t my_symbols socket memcpy strncmp lib_name symbol_count set_window_menu fill memmove fs_delete gui_draw_progress fs_rename free get_launch_args kernel_api_t sendto exec net_get_interface_info malloc memset mouse_cb_t fs_list process_events gui_draw_button tlen exit fs_create draw_image_scaled draw_image input_cb_t draw_text_clipped my_exports sprintf strchr cdl_main fs_read print uint32_t item_count menu_cb_t mem_total itoa dns_resolve paint_cb_t char strlen recvfrom strcpy draw_rect_rounded get_kbd_state bar_col realloc action_id GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection exec_with_args func_ptr long unsigned int draw_rect get_ticks pressed items get_fs_generation strcmp http_get percent strstr mem_used draw_text connect recv fs_write bind usr/lib/gui.c /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/lib usr/lib/../../sys cdl_defs.h    ���� |�  �              A�A�A�A�C0H<E@ADAHDLDPL0P<A@DDAHALAPF<E@BDAHALAPL<D@s0n
A�A�A�A�EOA�A�A�A� 8          <  A�BF���
�A�A�A�EX�A�A�A�         \            w            {                                             ��   t          �  ,           H                  ��!           7   x        @   w        V   {        l   h        �      <    �            �   \        gui.c sys my_exports my_symbols __x86.get_pc_thunk.si _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ gui_draw_progress gui_draw_button cdl_main  .symtab .strtab .shstrtab .text .gnu.hash .data .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                          �                 %         �  �  $                !   ���o   �  �  ,                +         �  �  �                   1         h  h                   :         t  t                    ?         x  x  �   	             H               @   	            P         @  @  ,                  X              �  �
                 d                �                 r              �   H                 �              "                     �              0"  `                 �      0       �#  Y                �      0       �(  g                 �              P)  $                 �   	      l  l                                t*  �               	              T+  �                                ,  �                  