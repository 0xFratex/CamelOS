ELF              �   4   �'      4    (                 �  �           �  �  �  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      VSR�   �à  �t$��   ��t0��������R��4$��   ���   ������T$ � ��[^��X[^��J   S  ��   ��t��j j j �t$,�t$,�t$,�P<��,�Ív �     �T$��   ��x���Ë$Ë$�[USR32] MsgBox:  
                                              A@(          ��V^�h��                    usr32                                 `                      msgbox                              create_window                   P   �                        �   ���o�      �     @  
   +            �                    ���o                                                           "   �               P        P   1      usr32_msgbox usr32_create_window cdl_main  H     �     �     �	       �  4           �       �  1   0  �   C   �   	P   U   o   o   o   o   o    int �  
�   �   �   o    n  �   �   �   o   o   o    �  �   �   �   o   o    	0�   �  �    �  #       1    #      #  1     	R  �  
R     4b  �  	o   �   b  1    �   r  1    �   #  	�	  �       -  �  F  j  V  �  \  �   p  �  !�  �  "�  �  %�     &�  $=  '�  (�   (�  ,T   )p  0�  *�  4R  +p  8U  .%  <x  /I  @8   0h  D�  1�  H�  2�  L�  3�  P�   4�  T(   5  X�  81  \�  9Q  `  :f  dy  ;�  hc  <�  l�  =�  pM   >�  tp   ?�  x   @Q  |5  A�  ��   B�  �  C  ��  F  �C  G  �E  H  ��  I<  �^   J  �  M�  ��  NZ  ��   Ox  �  Px  ��   Q�  �  R�  �o  S�  �i  T  �=  U,  �    VJ  ��   W�  �w   X�  �	  [\  �          C   &  &   +    C   F  C   &   2  V  C    K  [  o   p     a  o   �       u  �  �  o      �  o   �    �  o    �  o   �    C   o    �  o   �    o    �  8   %    o   o   E   v   �    �  I  o   o   o   o   o    *  h  o   o     o    N  �  o   o     o   o    m  �  o   o      �  �  o   o   o   o      �  �  o   o   o   o   o   o    �    8     o   �    r  �  1  C   o   &     K  C   K  &   P  6  f  �     V  �  �    &   k  o   �      &   �  �  �    o    �  �  �       �  o   �  �     �  &  �     �    o   �     &     7  7  7  7   o   "  o   Z  o   o   o    A  o   x  o   K  o    _  o   �  o   K  &  o   K  o    }  o   �  o   K  &  o    �  o   �  o   C   &  o   C   7   �  o     o   C   &  o    �  o   ,  o      o   J  �  �  �   1  �   ]}  	$_	{  �  _   �   _'C     \  _3Z  	,`	�  �  `     `)o    �   `6o   $#  `R�  ( {    `]�  �  O  sys �  �  {  �  1       �  `  B   �        �  �      �F	  
api '�  �  O  C   P   1   ��	  L  '  � 
w 2o   �
h 9o   � (      P   �L          
msg 2  �   I   :!;9I8   !I  'I  '   :!;9I  I  ! I/  	:!;9  
 :!;9I  $ >  4 :!;9I  %     $ >  & I  :;9   '  &       'I  4 :;9I  .?:;9'I@z  .?:;9'I@|   :;9I  .?:;9'@   :;9I�B                 C� LP�                   �           �     7   �          D   L   <   <   ^   7     !f	K) �: �= : f �0: V0<L�f<I>KJ,J�	� g net_get_interface_info memmove cdl_main set_window_menu draw_text my_exports strchr fs_delete get_fs_generation strstr http_get draw_rect_rounded fs_create win_handle_t kernel_api_t symbol_count sendto func_ptr paint_cb_t menu_def_t dns_resolve strlen bind itoa cdl_exports_t ping strcpy my_symbols long unsigned int close mem_used title fs_exists cdl_symbol_t recv mouse_cb_t strncpy get_kbd_state memset exec_with_args draw_image get_ticks realloc input_cb_t draw_text_clipped exec action_id get_launch_args item_count process_events items send char usr32_msgbox sprintf fs_list mem_total usr32_create_window strcmp free recvfrom draw_rect menu_cb_t print GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection memcpy exit socket uint32_t fs_rename lib_name fs_read label strncmp draw_image_scaled malloc connect version fs_write /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/lib/usr32.c usr/lib usr/lib/../../sys cdl_defs.h    ���� |�  <           P   A�A�A\G bA�A�B��AA�A�$       P   1   WBB B$D(D,D0F       �             �             �                                  ��	   �             ,        `  H                  ��#   �        ,   �         B   �         X   �        n   P   1     �   �        �       P      usr32.c sys my_exports my_symbols _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ usr32_create_window cdl_main usr32_msgbox  .symtab .strtab .shstrtab .text .rodata .gnu.hash .data .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                           �                  !      2   �   �                   -         �   �  $   	             )   ���o   �   �  ,   	             3               �                   9         �  �                   B         �  �                    G         �  �  �   
             P         @  @  @   
            X         �  �  +                  `              �  �	                 l              �  u                 z              �                    �                                   �              4  �                  �      0         (                �      0       /$  i                 �              �$  �                  �   	      �  �     	                           D%  �      
         	              &  �                                �&  �                  