ELF                4   �      4    (                 �E  �E           �P  �@  �@  �   �         Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      UWVS��L�  �Ð!  �$�|$d�t$l��4  ���   ��D  �$��(   �T$��<   1����
�T� �$��4  ���   ���D$��4  ���   =�� �  �����D$��$��D   �T$�D$������1���L$���C�<   ����D$���h&%%�VjPW�t$|�\$ ��4  �P@��4  �P@�\$ ��$   ���D$�8�%�U��-��� �O�L$(PjjPQ�t$|�ҋ�$�   �Y�� j��T$�����P�GPS�T$��4  �PD�T$��4  �@@���T$�:�X  �&%%���RjjP�W7R�t$|�Ѓ� j��T$�����P�GAPS�Ӌ�4  �PD�$�V�D$|��PPW�D$|��PP�\$ ��4  �P@��$�   �Z���$�   ��Z��h   ��F�PS�G
P�T$0R�D$ ��4  �P@��h333�jS����������P�t$0�D$ ��4  �P@�D$$� ���� ��u�l$�|$h�   �Q  �������,����)ݍF�D$�|7��t$1ۉ|$����D$�8�D$�ٸ������������)Ѝ Ѝ���)��D$����d~�d   �D$�ȸ��Q�������)ȋT$)�Ɂ�]+ ��i� ��QPURV�D$ ��4  �P@C�� ��<�m����$��4  ���   �D$�0����   �D$� ��;����D$�����\$(SP�ы|$��4  �@D���t$���uR�����h����R�t$$V�|$l�WdR�ЋD$��4  j�SV�D$|�   P�RD��l[^_]ý   �����   ������4$�����멋D$�u�����z �������  ���  �|$O$�D$����v�D$��8��w��$   �    Ð��$   �     Ív WVS�  �ƌ  �|$��4  1���D  ��D   f���    �    �
    @��<u��������j ������h�   h�  ��"���P�W<�� ������[^_�f��VS�t$��t&�D$�T$��f�@B9�t��8�t���)�[^Ð1�[^Ív UWVS����  ���  �t$0��tr�L$4��tj���t$<���  ���   ��Z�t$@���  ���   ��)�x=1��ŉ|$��v F�D$9�'�|$0�PU�t$<W�Q�������uމ����[^_]�f�1���[^_]ËD$�L$��u	�f�9�t
@���u�1�ÐS���  ��#  �D$���  ��uoǃ�     ���  ��������R���h@  j ���������  �P\��d  �     ��D  �     ǃ�      ���  ��3����T$ � ��[����t� ��t��d����T$��[��f���[Ív VSR�v  t  ��d  ���0�����  �t$�ҍ��  ��P�Qd����L$$�L� @���X[^�f�UWVS���  ��   �D$0�D$��d  ���~N���  �D$��1��
f�E��$9.~4���t$W���  �Pl����u��D� �T$�D� ��t��[^_]���v ��[^_]�S���  �ç  �T$�D$��dt@��etS��x9��  ��[�f������ ����D���  P�1�������[Ð����H���P��������[Ð����V���P��������[ÐVS�L$�t$�\$1����f��@9�t���u��� [^Ð�� [^�UWVS��@��  �  �D$�\$Tǀ�      h   j ���  �|$(W�ǋ��  �P\���; �5  ����b����|$$��h����D$(��  �D$�f��]�} �  ���t$,S�\$�z����Ń�����  ���t$0P���^�������t��p���  ����  �S���  �P����  �����D$�1��f�F@�T����t
��"t��u����߉\$ ؋L$� ���\$��o���PU������D$ �����M  9��4�����w����D$߉l$,�f��D$��8�   ���D$9��  ���t$ V�\$�����ƃ�����   9D$��   �D$��8�   ����   ����}���PV�R���������um���\$������PV�5����������p����P���e����D- �(���D$ ËD$�1���v ���?���@�T�T���.�����"u��$����P��t��\- ����D$ ËD$�1��@�T�T���b�����"�Y�����u��O����l$,�]�} �������<[^_]�1��n���U��WVS��L�H  ��N  �E��D  �M��    �8 ��  �������}��������M���d  �}���E�� �B	�z	 �b  ���u�P���������K  ���u�P����������4  �p��������PV����������  W��)��~�   �E�RV�}�W�q���Y^������R�E�P����������   ���u�P����������   �p��������PV�j���������   �Eċ ���(����U���W�����M��P���  �Pd���U���)�=�   ~��   �U�PV�Eċ �����M��D P�����XZ������PW���  �Pl�����U���������Eċ �����M��D P�������U�������e�[^_]�UWVS���  �ƈ  ��D  ���~N1�1ۍ�d  �D$�f�C��   9~1���t$8�D$�P���  �Pl����u׋D$�D ��[^_]Ív 1���[^_]�f�UWVS��   �  ��  ��$�   ������P���  ��4$���  ��������,$���  �_XV�|$W���  �Pd�<$���  ���   ����~�|�/t��������R�P���  �Pd�����  �pd��W���   ZY������R�P���$   ���  �P�ƃ�����   Ph   j V���  �P\��h�  VW���  �P ����~>� ��V�����4$���  �P���  �� ����$����   �Č   [^_]Ð��������P���  ��<$���  ��,$���  ����  �4$�P��1��Č   [^_]Ã����  ������R���1��܍v S���    �L$���  ��t#��t���  ��~������S���  PQ�RX����[�S�@  >  �\$�T$�L$���  ��t�@L��t�\$�L$�T$[���[�f�S�    �\$�T$�L$���  ��t�@L��t�\$�L$�T$[���[�f�UWVS��8�  ���  ������P���  ����  ������  ��D  �|$Ǉ�      ��h   �P�ƃ����g  Ph   j V���  �P\��j@V�G(P���  �P(������  �D$    ���  ������|$������|$�t$�T$f��> ��   ���t$V�Pl������   �~0�����  ��u7���t$�L$���   U�Pl�����  ���  �L$���    ��   �L$���  ��?F�i�T$���  ��V�,	����T$���   Q�Pd�T$Չ�$  �F(��(  �����  �D$�T$��@9T$�.����t$��V�P�D$ǀ�   ����ǀ�       ���  �������$�����,[^_]Ív ��V���   �D$,�,$���  ���   ��9D$�y�����U�L$()��P���  �Pl�����W������  ���������  �_����VS���  �Î  ���  �����R������  h   j ��D  V�P\�    ���  ��*����$���[^�f�UWVS���2  ��4  �D$ �l$$�|$(��D  �   �C    ���  �Rd��tb��P�CP�ҋ��  �@d����tX��U�S(R�Ћ��  �@d����t6��W���   R�ЋD$<���   ƃ�    ���������[^_]Ð��B���떍������G����VSQ�z
  �À  �t$�t$ �t$ �t$�t$�!�����D  �@   ����t���  �t$�   �D$�BdZ[^��f�X[^�UWVS���&
  ��   ������S��D  �n(U���  �Pl����t=��U���  ���   ����~-�P��|'/u�E�Ht)�T(��/u��D( ���������[^_]�u�V)�����u���S�F(P���  �Pd����f��D' ��1�븐WVS�v	  ��|  ����D  �~(W���  ���   ����~ �|'/t��������R�P���  �Pd�����  �xd����(V���   ZY�t$�V���D�����[^_ÐUWVS��   ��  ���  ��D  ���   ��x;��  �  ���C(P�l$U���  �Pd�,$���  ���   �ǃ����  �|/t6��������R�T$U���  �Pl����t���T$R�W���  �Pd���{��tb�����   W���  ���   ����t7���  �pd��U���   ZYW�P�֋��   ����t	��U�Ѓ��    �Ĝ   [^_]Ív ���   ��x�;��  }����  �pd��U���   ��XY�?������   P�R�f�� �����$  ������������   P���������f��!�����������PU���  �Pd���{�������c����v UWVS��,�N  ��T  �|$@�t$D��D  �E ���C  ���  ���[  �L$H��p������T$����L$�T$L���������1�T$��jh   @h,  h�  �LQ�L$ �TR�PT��jh����h,  h�  �t$,V�|$$W���  �RT��h����jh�  VW���  �R@��h����jh�  ��,  RW���  �R@��h����h,  jVW���  �R@��h����h,  jV���  R���  �R@�|$(��
��jh����jj�V
RW���  �RT�t$4���� h   ���R���RV�D$�PR���  �RDh   ��URV�D$$�P2R���  �RD��h�   hfff��U(RV�D$$���   R���  �RH�t$4��(�� �}��  �D$
   ��   ��j�P�D$h|  VW���  �R@��h����jh|  VW���  �R@��h����jh|  �D$�PW���  �R@�D$4��*�� 1���]����L$��O����L$�|$���g�v �L$�D$��jjW�D$�PRQj ������ h   ��D$������   P�GP�D$��#P���  �PD�D$�D$�����L$9�td�t$��   9��  ~R9��   u'��h�׳�jhz  �G�P�D$$��P���  �P@�� �6�0����$  ���C����L$�>���f��D$��  �}��   �L$�D$���   h   ���T���RW�t$�VR���  �RD�D$$�   �t$��<�$����jh�   P�D$ V���  �R@��h   �jh�   �D$PV���  �R@�� h   ����   RW�t$�VAR���  �RD���L$��jh����jj<Q�L$ �|$$���   R���  �RT�t$4��  �� h   ���Z���RV��  R���  �RDXZjh�z �jj<�L$Q��@  R���  �RT���  �RD�� �}t<��B���j�PV�D$O  P�҃��   ��,[^_]�f��D$   ��   �G���f���M�����1���,[^_]�f��  �»  ��D  � ��t1����  ����Ív UWVS���  �Ì  �T$8��D  ���tg�D$0-�  ��9�S���  9�|I�|$4��,  ��;|$<7��,  ;t$<|+�p	9���   �p(9�|)�w	;t$<} �w;t$<|�����f��   ��[^_]Ív �q�t$N�
  ��   ��|  9�|�o(9l$<|v�;t$<|n�T$<)�����������   x�9��  ~�9��   ��   ���   �|$u�k�0��$   �x���PP���  ���   R���   R�Pd���V���f���  ���   9�},��6  9�|"9t$<�0�����  ;l$<|�    �������?  9��
���|  9������9t$<�������  ;|$<������������������   �����k�0��$   u�|$ �>����у����   P�4���������S���   �§  ��D  ���t�|$tn�|$
t�{t�   ��[Ív ���e�����v �����  ���   R���   ���|$t0�L$�Q���^w���>��L$���   Ƅ�    �f��    뗅�~�Ƅ�    뉋$Ë$Ë4$Ë$Ë<$�  CPU % MB Used CPU RAM Activity Monitor [FW] cm_init: Done.
 fs_new_folder fs_new_file <Menu name=" </Menu> <Item label=" id=" <key> </key> <string> </string> CamelMenuDef [FW] Loading config for:  / Info.clist [FW] Picker Refresh...
 [FW] Picker Refresh Done.
 . * [FW] Dialog Init...
 [FW] Dialog Init Done.
 Open /home Save ^ Name: Cancel    [FW] WARNING: cm_init called twice!
    [FW] cm_init: Setting up framework...
  [FW] Failed to allocate config buffer
  [FW] Config not found (or empty):   [FW] Config loaded successfully.
   %   '   !                                                   &                $           %      	      #                                                                                                                 
          "                                                      %             %� �-&�C @  1+�  H                           
                                                                                      "   &           2�?���!wp���Lʽ|����h#�bϐtz5ӝ���rMw9J/q|aI�b*�|EI�%+R�E���P�Y�^47(2ӏigswї|)��� c��Wm+�c%1hjі����"Sn7���K��	9�xy�U	��Bd8��J��|iB����            Waterhole                                  �   :      �  �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �  ���o�     |C     A  
              �E                     ���o                                                           �   �  �    ^    :  @    �    {     �   x  8            �    �  �  %        1   	    o  \  �     B   �  �     �  �  �     f    :       D  �  3    �  <  �    .  �  :     &   �  E     
   �"  �     �   p  |     V  �#       `    V     �      N        �!       V   p  �     L   P       �  �  �    �   �  �     �     v     /     u         D     ~    \     �   �  �    �    �    �  p  �        �!  �     �   @
  �       X  :     !   �!       8   �  5     s   �0        on_paint cpu_hist head ram_hist mode on_mouse cdl_main my_memcmp my_strstr my_strchr cm_init actions action_count config_count cm_bind_action execute_action_by_id internal_menu_callback strncpy_safe parse_menus_from_string parse_plist_xml cm_get_config cm_load_app_config cm_apply_menus cm_draw_image cm_draw_image_clipped cm_picker_refresh cm_picker cm_dialog_init cm_dialog_open cm_dialog_save cm_dialog_up_dir cm_dialog_select_dir cm_dialog_submit cm_dialog_render cm_dialog_handle_mouse cm_dialog_click cm_dialog_input �!     �!     �!     �!     ~       d             }      �  1   �  Q   C     	P   U   o   o   o   o   o    int �  
�   �   �   o    =  �   �   �   o   o   o    �  �   �   �   o   o    0�   K   �    Z  #   	    
1    8    	  #  
1     	R  �   
R   �  4b  �  	o   � 	  b  
1    	�   r  
1    )   #  �	  �     /  -  R  F  �   V  h  \     p  �  !�  �   "�  �  %�   	  &�  $H  '�  (m  (�  ,�   )p  0�   *�  4A   +p  8^   .%  <�  /I  @�  0h  D�  1�  H�	  2�  Lw  3�  P2  4�  T�   5  X6  81  \�   9Q  `+  :f  d   ;�  h�  <�  l�   =�  pl  >�  t�  ?�  x�   @Q  |�  A�  �  B�  ��  C  ��  F  ��  G  ��  H  �D  I<  ��  J  �    M�  �z   NZ  �  Ox  ��  Px  �  Q�  �<   R�  �"  S�  ��  T  �   U,  �  VJ  ��  W�  ��  X�  �P  [\  �          C   &  &   �    C   F  C   &   2  V  C    K  [  o   p     a  o   �       u  �  �  o      �  o   �    �  o    �  o   �    C   o    �  o   �    o    �  8   %    o   o   E   v   �    �  I  o   o   o   o   o    *  h  o   o     o    N  �  o   o     o   o    m  �  o   o      �  �  o   o   o   o      �  �  o   o   o   o   o   o    �    8     o   �    r  �  1  C   o   &     K  C   K  &   P  6  f  �     V  �  �    &   k  o   �      &   �  �  �    o    �  �  �       �  o   �  �     �  &  �     �    o   �     &     7  7  7  7   o   "  o   Z  o   o   o    A  o   x  o   K  o    _  o   �  o   K  &  o   K  o    }  o   �  o   K  &  o    �  o   �  o   C   &  o   C   7   �  o     o   C   &  o    �  o   ,  o      o   J  �  �  �   1  �   ]}  $_	{  �   _   �  _'C        _3Z  ,`	�  �   `   4   `)o    �   `6o   $  `R�  ( {  l   `]�  �  O  sys �  �#  	o   �  
1   ;    �  �"     �  �!  �   o   �!  �   o   �!  �   P�  `!  �  Q�    u   ��	  api Q'�  � win TC       +   i So           !_  I�	  x o   y o   btn !o    "�      �  �   x o   � y o   �w !o   �h (o   ��  &   $       �  &   8   2   �  	o   Y   U   mx (	o   v   l   mw )	o   �   �     1
7  �   �   �   2	o       buf C
  �@   i 5o   K  E     idx 6o   d  b  val 7o   �  |  �  :o   �  �  bx ;o   �  �  by <o   �  �  col >&      #�	  �  E   ��	  � �	  ��	  �$�	  �   '   I�	  �  �  �	  
    �	         �   �  4d  t      �    �  �  2   �  Q   E   5  	S   X   r   r   r   r   r    6int �  
�   �   �   r    =  �   �   �   r   r   r    �  �   �   �   r   r    0   K       Z  #   
    2    8  7  
  ,  2     ]  �   
]   �  4m  �  	r   � 
  m  2    
�   }  2    )   ,  �	D  �  T   /  o  R  �  �   �  h  �     �  �  !�  �   "�  �  %   	  &  $H  '!  (m  (:  ,�   )�  0�   *�  4A   +�  8^   .g  <�  /�  @�  0�  D�  1�  H�	  2�  Lw  3  P2  45  T�   5Y  X6  8s  \�   9�  `+  :�  d   ;�  h�  <�  l�   =�  pl  >�  t�  ?  x�   @�  |�  A,  �  B@  ��  CU  ��  F_  ��  G_  ��  H_  �D  I~  ��  J_  �    M  �z   N�  �  O�  ��  P�  �  Q�  �<   R
  �"  S7  ��  TZ  �   Un  �  V�  ��  W  ��  X  �P  [�  � O  O     D  E   h  h   �  Y  E   �  E   h   t  �  E    �  8�  r   �  O   �  r   �  O  O   �  �  �  r      �  r     O  �  r    �  r   !  O  E   r      r   :  O  r    &  9   g  O  r   r   G   y   �    ?  �  r   r   r   r   r    l  �  r   r   O  r    �  �  r   r   O  r   r    �  �  r   r   O   �    r   r   r   r   O   �  5  r   r   r   r   r   r      T  9   T  r   �    }  :  s  E   r   h   ^  �  E   �  h   �  9x  �  �  O   �  �  �  O  h   �  r   �  O  O  h   �  �  �  O  r    �  �    O  O   �  r   ,  �  O  :   h  @  O   1  U  r   �   E  ;&   Z  y  y  y  y   r   d  r   �  r   r   r    �  r   �  r   �  r    �  r   �  r   �  h  r   �  r    �  r   
  r   �  h  r    �  r   7  r   E   h  r   E   y     r   Z  r   E   h  r    <  r   n  r    _  r   �  �  �  �   s  �   ]�  �  �  T  0-�  �   .�   =  /r   (�  0r   , 
  �  2   '  �	    	r    �   	r   �  
  L  
�	  (�	   
�	  �R	  !
�	  ��  $	r   �0  %	r   ��	  (�  ��  1�	  �<g  2	r   � 
  �	  2    
  �	  2   ? 
  �	  2    
�  �	  2   ?   3�  =�  6�	  /  �  �  1  K  �  �  &   >sys �  �@  $2	I
  &id 3  �  4�    ^  5)
  
I
  e
  2    �	  7U
   :  �  8r    :  
}  �
  2    S  :�
  �<  -  ;r   d<   >�
  &key ?  �  @
�
    
  �
  2   � _  A�
  
�
    2    �  C�
   1  ?  Dr   �0  ?�	  O�#      �r   �  �   ��  key �r   � �   }  len �r   @  <   /  �    �  fr     �  ��  	?	  fr   � 	4	  f$r   �mx f/r   �my f7r   �x i	r   a  O  y j	r   �  �  (  u	r         v	r   ;  5  fy �	r   W  U  �   }  idx zr   c  _  �  {r   �  �  �  �  �  �   !�  &  �   i�  �  �  �   !�  1  �   j�  �  �  �   �  #   @�  Er   �  %   �  mx E r   � my E(r   �btn E0r   �  �  �r   <  �  ��  	�	  �r   � 	E	  �%r   �	?	  �0r   �	4	  �;r   �x �	r   �  �  y �	r   G  ?  (  	r   �      	r   �  �  D  	r   �  �  A�  	r   fy 0	r   �  �  "a  �   S  i r       �   idx r   8  4  iy  r   S  G    (O  �  �  �  ^    !�  u  �   �v  �  �  �   '�  �  �   ��  �  �    (�  ��  �  ��  �  �
�	  ��~len �	r   �  �    �   #s  �  {   �#  	  �'O  � len �	r   �  �  B�  w �     C�  �=  )len �r    DX  �  \   ��  �  �!O  �  �  �  �4O  �  �  	�  �KO  �	K	  �eO  �cb �~�  �;  �   #=  �\  �   �  	�  �!O  � 	�  �4O  �	K	  �KO  �cb �d�  ��     E�  �  V   �(  [�  3  ��  F@d�  �  e�   �  f&   (�  g&   ,�  h�	  0*uid i�	  1�  j�	  2*gid k�	  3�  l�  4 G	  m4    o	r       "	  p�  .  $  �  F  u	r   `  T     i wr   �  �  �   =  {r   �  �  �  �r   �  �  �   i  �  �r   �  �  :	  �r   
       F   idx �r           
&   �  2    +	  H�  :   �^  U  H&
       �   H8O  ;  1  x HBr   h  b  y HIr   �    dw HPr   �dh HXr   �cx H`r   �cy Hhr   �cw Hpr   � ch Hxr   �$,�  -��  +�	  EX  :   ��  "	  E
  �  �  �   E2O  �  �  x E<r   �  �  y ECr   �  �  	�  EJr   �	�  EUr   �,�  -��  #�  "  D   �  	)	  "E   �  $�  �r   �  �  �o  �	  �$O  V;  
�	  ��~)len r   V  
�  V�  	r   P $  �O    v   ��  key �'O  �   O   i �r     
    %  ��  �  �2  xml �$�  � ptr ��  &    I   �  ��  O  E  {  ��  z  t  Y     �	  �r   �  �  i �r   �  �  �  ��  �  �  m	  ��  �  �  i     	  ��  	  �  �  �r   $	   	  �  ��  ?	  3	  �  ��  �	  |	  "�	  H   �  k �r   �	  �	   "�	  L   �  k �r   �	  �	   +	  �  f	  �  �	  �   �  �   >  �  Z  �    %F  �@
  �  �j  buf ��  �	  �	  ptr ��  �	  �	  t   �  ��  
  
  m  ��  
  
    ��  !
  
  v	  �  �@Z  �r   -
  )
  s  ��  R
  P
  �  ��  `
  Z
  ]	  ��  z
  v
  �  �r   �
  �
  �
  �  �
  �  �
  �    j    �  0  �  N  �  �  j  �  �    H�  �x  8   ��  I�  ��  �
  �
  src �+O      n �4r   F  <  i �	r   s  m   J�	  m�  .�  m!r   .�	  m/r   Kid }O   /l  cp  |   �2  id c'O  � >   i dr   �  �    %,  \   N   �c  Z  \!O  � �  \3�  � /%  Hp  �   ��  api H�  �  �  �  Ir   `<   0i  &�  P     ��  s &O  �  �  c &$r   �  �   $�  �  �  �   �X  �  O  � L  3O  �'  	r   �  �  �  	r   �  �     8   i  r       /  X    0_  r   �  5   ��  s1 �  � s2 +�  �n =h  �p1 O      p2 O  '  %  �  &   i h  6  .    L�	  r   �  Mval !r    N�  �  �   �z  1�  � 1�  �2�  f  `  O�  `   `     mg  �  �  �  �  �  �  3�  o  �   ?  �  W  �   P#  p  �   �31  '#  �   �   ��   21  �  �  �         I   :!;9I8   !I  'I  '   :!;9I  4 :!;9I�B  4 :!;9I�B  	I  
! I/   :!;9I  :!;9  4 :!;9!I?  $ >   :!;!� 9I   1   1�B  4 :!;9I  4 :!;9I  U  %     $ >  & I  :;9   '  &       'I  4 :;9I  .?:;9'I@|     !.?:;9'   ".?:;9'@|  #.1@z  $1R�BUXYW    I   :;9I8   !I  H }  'I  '  4 :!;9I�B  4 :!;9I�B  	 :!;9I  
I  ! I/   :!;9I  4 :!;9I�B   :;9I  4 :!;9I�B  $ >  U   1�B   :!;9I�B   :!;9I8   :!;9I   :!;9I�B  U   :!;9I  :;9  4 :!;9I?  4 :!;9I  4 :!;9I     :!;9I�B  :;9!	   .?:!;9!'I@|  !1R�BUX!YW  "  #.?:!;9!'@|  $.?:!;9'I@|  %.?:!;9!'@|  & :!;9!
I8!   '1R�BUX!YW  (.?:!;9!@|  )4 :!;9!	I  * :!;9!I8  +.?:!;9!'@z  ,H}�  -I ~  . :!;9I  /.?:!;9!'@  0.?:!;9'I@z  1 1  24 1�B  34 1  4%  5   6$ >  7& I  8 '  9&   :   ; 'I  < :;9I8  =4 :;9I?<  >4 :;9I  ?4 G:;9  @.?:;9'I@z  A4 :;9I  BH }�  C.?:;9   D.?:;9'@  E. ?:;9@|  F:;9  G :;9I  H.?:;9'@z  I :;9I�B  J.?:;9'   K4 :;9I  L.:;9'I   M :;9I  N.1@z  O1R�BXYW  P.1@|   ,           ��0���P     djPj���       p�p D%���Q��p D%�    ��P���P�          ��� #P���P������� #P���� #P�          ���P���P�������P����P�     ��������          ��s <���
�d<���U��s <���U      ��0���S��S  ���!  s "<�  ���!  s "<2$��"��$�!  s "<2$��"d-( �     ��P����  ��V   ��R    ��� ���     ������     ������ �
            �/�/P�0�0P                   �+�,P�,�,
� 
�1&��,�,P�,�-
� 
�1&��-�.P�.�.p�}��.�.
� 
�1&��.�.P�.�.
� 
�1&�        �+�+
�
,1&��+�+w 1&��+�,
�
,1&��,�.
�
,1&�    �,�-�
,1&#(��.�.�
,1&#(�      �,�,ȟ�,�,V�.�.ȟ   �-�.V    �,�-	�u D��.�.	�u D�         �,�,
r �$  "��,�-R�-�-�$  �.�.R    �+�+� 
���+�+P �+�+�
,�             �"�"Q�"�#�H�#�%�D� "��%�*�
�1&� "��*�*�D� "��*�*�
�1&� "�         �"�"R�"�$�T�$�*�
,1&�"��*�*�
,1&�"�         �$�&V�&�*�T#(��*�*V�*�*�T#(�    �$�%ȟ�*�*ȟ    �%�*D��*�*D�         �'�(Q�(�)�L�)�*�T#���*�*�T#��        �%�&0��&�&�D�&�&P�&�(�D     �&�&V�&�(V            �&�&w~��&�&wj��'�'w~��'�'P�'�'���'�'w~�   �&�&Q �!�!�
�� �"�"�
,�         ��P��W�!�!P�!�!W   ��P     ��� ���      ������    ��@���@�         ��P��V���X���X��V             ��P��R���L���L��P��R          ��0����D��R���D��0�       ��w 1���W��W    ��0���0�     ��P���\   ��P   ��Q     ��� ���            �����S�����S���       �����R��R     �����Q     ��� ���            �����S�����S���       �����R��R     �����Q    ��0���S        ��S��S������S           ��U��P��U���\��U       ��P��V��V       ��S��	d<  1���S      ��0���P��0�     ��P���@     ��V�	�	V         ��	V�	�	v{��	�	P�	�V     ��	U�	�U          �	�	P�
�
P�
�
p��
�
q��
�
q p "#��
�q p "#�        �
�
P�
�
p��
�
q��
�
q p "#��
�
q p "#�    �
�
0��
�P    �
�
0��
�
P   ���     ��P��P   ��P     ��P��V   ��P  ��p v ���p v O-( �   ��P       ��V��P��V     ��P��R       ��p v ���r v ���u�v �-( ���r v �-( �           ��� ��Q��� ��Q���            �����V�����V���           �����S�����S���      ��0���P��P    ��0���U       ��� ��� ���      ��� ��P     �����Q     ozPz�W     ��P��U    ��0���V  5�   5�      0�p � �	p � #�*p � �      ��p 0r 8$"�<  "���p 0� 8$"�<  "����0� 8$"�<  "�   ��R���  ��e�           ��P��p���P��P��P��R��P                  }              �       �            .         ���� ������ ���� �         ���� ������ ������ ��	�	� ���� ���� ���� ���� ���� �!�!�!�" �"�"�"�" �%�&�&�' �+�+�+�+ �+�+�+�+ �,�-�.�.�.�. �/�/�0�0 �    7   �         M   V   	   	   i   +     � �( J. �u �ufg �>f�#�JJ=<
�i�,�� < ./,� � X!�	�u	,J>�?7 ��?(� tK	��1	 vy�/�	rf��t		h/	J�� v   .��% �/ � < t tK� � fK�t l  e� -� � `�&%��s	t	Yt X$  � +$ 	�,O!	g	 # �. 2 �=  t  Y�K =
 �    <   �         �   �   |   |   i   �   @ �  g	 "     	Y.< J& * <1I/;h! ��K�g	  X.! �  	�f � �t& yX5'��	�	K
 s4!./��	h�����f�/I	r. J . J� qJJ@���Y<f&J�K .�g+h�	 t# f  	u u�" J" p X9�i]^ J�r;<X��	sf�<nf	
�D7k� ' �/ # <   J <+ J/=  	-.=  )7 ���x'��	!<P	��X	/	�	�u>!f�(�11<-h8) - 1I1. J1 X['<�<K��fN�-�<h�"/ ��Ju�!{Y�: $ : < � : t�CG : I$ : J* � �w< $ < < �K?C < I$ < J+ �< � �	J<P2�Y�!�tg�#%1�
�	[<S	�	�	�#	�  �1 	>!	�	�K	��.	�	�#	� �0 	?!	!	�<.�1J��y<z�2. i .�A<  ,;�!	 �# �  	�&tf �7 t> �Js/5��. �K �� f. tv� ��!�"/{L��f��	s�;  S �	�	fgx<.	l�<	f�'�!	f JKf	KL\Xgf J <  J J JK  = |=gf J <  J J JK  = <!�	f�@)��"L	 ���	t<	� �	�2	zd<0 J�= b  �Y,�/J.K+�)� cf J J !v��f�j���g�?Jf< � � � ff�f�<fgf�h���u� J�� t�� t��!uu z� � ���!K� t  f J �= ;KL!	 �s�- � <9 �   + . J
Z%Zu }+ .g J t	�&	Y &-.0<�� t9 t ��)� ��Y�L�' J�K �/ t J, <	u��	| Xu%� � yf/f% t�
f	s�f+ J�%� �h. �	m�8��M<t�t	g��<B��� � f��|��|�	 �.��|��|�	 �.x�M'����J�J$�&	u	I[����
 �E . � J	�w:�	�) pX J J <	�	�	���@X�	@2E� � �	�	���#��('*"� � f���0 O� .�+ ��� .5��� J�;OY�L�{��{�.��{� J fH�{�." �6 f, fi< � <( J" <: f0 <	gYF );XN�t	s[$  f	F( @G f8 .	gfX	[f .��*iS t4 <�.Vft��	if2 J f7 JO �C f	g	gjf1 � X6 �N �B f9 c� �0 s
�0<��E<tf'���LyyxfX	p�u	]<f	��t, XY-�-�	p	g. J: 
 ping close ram_hist strncpy cdl_symbol_t menu_def_t version send fs_exists label win_handle_t create_window cdl_exports_t socket memcpy mode strncmp lib_name bar_w symbol_count set_window_menu head memmove fs_delete exports fs_rename free get_launch_args kernel_api_t sendto exec net_get_interface_info malloc memset mouse_cb_t fs_list process_events on_mouse exit fs_create draw_image_scaled sb_w input_cb_t draw_text_clipped sprintf cdl_main fs_read print uint32_t item_count menu_cb_t mem_total itoa dns_resolve data paint_cb_t symbols strlen recvfrom strcpy draw_rect_rounded get_kbd_state realloc action_id GNU C17 13.3.0 -m32 -march=i386 -mtune=i386 -mno-sse -mno-sse2 -mno-sse3 -mno-ssse3 -mno-sse4 -mno-sse4.1 -mno-sse4.2 -mno-avx -mno-avx2 -mno-mmx -mno-3dnow -mno-80387 -msoft-float -mno-fp-ret-in-387 -mgeneral-regs-only -minline-all-stringops -g -O2 -fno-stack-protector -fno-builtin -fPIC -fno-tree-loop-distribute-patterns -fno-strict-aliasing -ffreestanding -fno-asynchronous-unwind-tables -fno-exceptions -fno-unwind-tables -fomit-frame-pointer -fno-tree-vectorize -fno-tree-loop-vectorize -fno-tree-slp-vectorize -fstack-clash-protection exec_with_args func_ptr draw_rect get_ticks get_fs_generation bar_h strcmp on_paint http_get mem_used draw_text connect recv cpu_hist fs_write bind key_content_end hlen cm_bind_action clist_path parse_plist_xml file_buf my_memcmp my_strchr cm_dialog_select_dir file_picker_cb_t perm visible_items start_dir long long int cm_dialog_submit show long long unsigned int dates my_strstr parse_menus_from_string active cm_dialog_input selected_index config_count current_dir cm_dialog_save entry_count val_tag name_ptr full_path value attr initialized real_idx nlen default_name menu_end key_tag size short unsigned int i_idx cm_dialog_handle_mouse dirname max_read file_picker_t cm_init temp_menu_count cm_dialog_open needle temp_menus action_bind_t execute_action_by_id entries strncpy_safe cm_dialog_click filename title id_p req_h haystack dest menu_idx cm_picker menu_tag req_w cm_dialog_up_dir cm_get_config list_h cm_picker_refresh list_y unsigned char is_dir item_h short int buff klen config_pair_t key_content_start icon lbl_p scroll_offset action_count cm_dialog_render cm_dialog_init cm_apply_menus func val_content_start vlen cm_load_app_config item_tag cm_draw_image_clipped buffer win_handle win_h flen win_w win_y filter filter_ext val_content_end item_ptr key_name raw_entry_t internal_menu_callback filename_input app_bundle_path win_x cm_draw_image item_idx actions safe_div2 usr/apps/waterhole_cdl.c /home/gustavo/Documentos/AIProjects/camelos/CamelOS usr/apps usr/apps/../../sys cdl_defs.h usr/lib/camel_framework.c usr/lib usr/lib/../../sys camel_framework.h       ���� |�            �  A�A�A�A�C`�lEpAtBxA|D�cl[pBtBxA|D�O`BdKhDlAp]`UlApBtBxD|D�E`BdKhDlApStHxA|H�dlEpDtAxD|E�PlEpBtAxN|D�X`�lApAtAxA|A�S`|hElApR`UdAhElHpNtAxA|J�FA�A�A�A�A`����         �  E   @         u   A�A�A�CFB F$E(E,G0FG�A�A�       �            �            �        ���� |�  ,   �  �  5   A�A�k
�A�BC�A�   l   �  �  �   A�A�A�A�C0^<D@O<D@O0a4A8D<A@H0K
A�A�A�A�CGA�A�A�A�     �  P     D   �  p  �   A�ClG EEBF @A�B�W
A�DCA�0   �     N   A�A�AZJM VAA�A�X   �  p  |   A�A�A�A�C0|8D<A@L0W
A�A�A�A�ECA�A�A�A�T   �  �  �   A�Cl
A�CCW HC
A�BCG HC
A�BCG HCA�,   �  x  8   A�A�k
�A�BF�A�   �   �  �  �  A�A�A�A�CTaXB\K`NP}XD\A`NPKXD\A`JPgXK\A`LPAXD\A`NPiXG\A`JPGXK\A`JP�
A�A�A�A�A(   �  @
  �  A�BF�����A�A�A�X   �    v   A�A�A�A�C0w8D<G@L0O
A�A�A�A�DEA�A�A�A��   �  �  �  A�A�A�A�F�Y�e�A�A�E�Z�N�G�C�K�L�A�G�A�G�C�W�I�E�B�A�L�E�A�A�L�K�A�e�K
A�A�A�A�BC�G�m�H
A�A�A�A�AC�M�E�,   �    D   A�ClAGA FCA�     �  X  :   A�t
�CA�   �  �  :   A�t
�CA��   �  �  3  A�A�A�A�CLRPQ@_LEPH@IDEHBLAPLDBHALDPN@@HDLAPF@]HDLKPF@~HALTP[@bLAPo@C
A�A�A�A�DCLAP\@MHALJPL@  4   �    V   A�A�CX EKBG ]A�A� d   �  \  �   A�A�A�A�C z(A,D0N G(A,D0N G(A,G0]A�A�A�A�B ����  D   �    \   A�A�ASDDD U[
A�A�DAA�A�   X   �  p  �   A�A�A�A�C(R,J0L G,A0O m
A�A�A�A�AO(A,D0L  T   �    {   A�A�A�NJ ONGC LLD GADC JA�A�A�   �   �  �  �  A�A�A�A�F�j�D�E�]�R�G�E�L�G�E�C�L�J�G�O�P�A�G�A�A�C�K�G�A�E�L
A�A�A�A�D^
�A�I�A�P�C�DZ�H�J�M�G�A�L�     �  <  �  A�A�A�A�C@`HBLEPETEXE\I`FHBLEPETEXE\E`LLEPBTEXA\A`LLEPBTEXG\A`LLEPETBXA\A`LLEPETBXA\G`SHBLEPBTBXD\A`S@EDGHALHPNTDXA\H`LLEPETDXA\K`S@ZLBPATIXA\A`LLEPBTEXA\A`LLEPBTEXG\A`S@lHBLBPATHXA\B`H@EDQHDLHPW@eLEPBTEXD\H`L@JDGHALHPbTEXA\E`LLEPBTEXE\A`L@EDGHALHPL@GHBLEPBTBXA\O`V@EDGHALGPJLAHBLEPBTBXE\G`U@NDAHALJPE@H
A�A�A�A�CaA�A�A�A�   �  �  %   T   �    �  A�A�A�A�C0�
A�A�A�A�Dy4A8N<G@F0�<H@H0(   �  �  �   A�Cs
A�DOM I    �  �        �  �        �  �        �  �        �  �                                 ��   �#          `!  ,                 ��   �@       /   `<       =   d<       M   �<                    ��X   �        n   �        �   �@       	 �   �        �   �        �   �        �   �!        �   @
  �    �   �  �       <  �       :       #  �  %     :     N     I  x  8     V  �0       c  P       m  �  3      X  :     �  �  �    �    \     �  p  �     �  �  �    �  �  E     �  \  �     �  �!       �  �!       �  �  :       �"  �       p  �         v     -    �    =   :  @    E  �  �     O  p  |     d  �  �    w  �#       �      �    l   1   	    �    u     �  �!  �     �    V     �    D     �    {     �  �  5     �  �  �      waterhole_cdl.c sys exports camel_framework.c initialized.0 temp_menu_count temp_menus __x86.get_pc_thunk.si __x86.get_pc_thunk.di _DYNAMIC __x86.get_pc_thunk.ax __x86.get_pc_thunk.dx __x86.get_pc_thunk.bx _GLOBAL_OFFSET_TABLE_ parse_plist_xml cm_dialog_input cm_dialog_render action_count cm_dialog_handle_mouse cm_bind_action strncpy_safe config_count my_strchr cm_picker_refresh cm_draw_image cm_dialog_submit cm_dialog_save cm_init parse_menus_from_string on_mouse cm_dialog_open mode head cm_draw_image_clipped cpu_hist cm_dialog_up_dir cm_get_config cm_dialog_click actions my_strstr execute_action_by_id cm_load_app_config cm_picker on_paint cdl_main ram_hist cm_dialog_init cm_apply_menus cm_dialog_select_dir my_memcmp internal_menu_callback  .symtab .strtab .shstrtab .text .rodata .gnu.hash .data .got .got.plt .bss .dynamic .dynsym .dynstr .debug_info .debug_abbrev .debug_loclists .debug_aranges .debug_rnglists .debug_line .debug_str .debug_line_str .debug_frame .rel.dyn                                                          �                 !      2   �  �,                  -         �  �.  8  
             )   ���o   �  �/  \  
             3         `!  `1  ,                   9         �!  �1                   >         �!  �1                   G         �!  �1  �                  L         �@  �P  �                U         A  Q  p              ]         |C  |S                   e              �U  @%                 q              �z  0                               �                   �              )�  @                  �              i�  �                  �              f�  e                 �      0       ˣ  �	                �      0       ��  �                 �              x�  L                 �   	      �E  �U      
                           ĺ  p              	              4�  �                               $�  �                  